// megafunction wizard: %ALT2GXB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt2gxb 

// ============================================================
// File Name: altpcie_serdes_2sgx_x1d_10000.v
// Megafunction Name(s):
// 			alt2gxb
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.1 Build 198 11/07/2006 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcie_serdes_2sgx_x1d_10000 (
	cal_blk_clk,
	fixedclk,
	gxb_powerdown,
	pipe8b10binvpolarity,
	pll_inclk,
	powerdn,
	reconfig_clk,
	reconfig_togxb,
	rx_analogreset,
	rx_cruclk,
	rx_datain,
	rx_digitalreset,
	tx_ctrlenable,
	tx_datain,
	tx_detectrxloop,
	tx_digitalreset,
	tx_forcedispcompliance,
	tx_forceelecidle,
	pipedatavalid,
	pipeelecidle,
	pipephydonestatus,
	pipestatus,
	pll_locked,
	reconfig_fromgxb,
	rx_ctrldetect,
	rx_dataout,
	rx_freqlocked,
	rx_patterndetect,
	rx_pll_locked,
	rx_syncstatus,
	tx_clkout,
	tx_dataout);

	input	  cal_blk_clk;
	input	  fixedclk;
	input	[0:0]  gxb_powerdown;
	input	[0:0]  pipe8b10binvpolarity;
	input	  pll_inclk;
	input	[1:0]  powerdn;
	input	  reconfig_clk;
	input	[2:0]  reconfig_togxb;
	input	[0:0]  rx_analogreset;
	input	[0:0]  rx_cruclk;
	input	[0:0]  rx_datain;
	input	[0:0]  rx_digitalreset;
	input	[1:0]  tx_ctrlenable;
	input	[15:0]  tx_datain;
	input	[0:0]  tx_detectrxloop;
	input	[0:0]  tx_digitalreset;
	input	[0:0]  tx_forcedispcompliance;
	input	[0:0]  tx_forceelecidle;
	output	[0:0]  pipedatavalid;
	output	[0:0]  pipeelecidle;
	output	[0:0]  pipephydonestatus;
	output	[2:0]  pipestatus;
	output	[0:0]  pll_locked;
	output	[0:0]  reconfig_fromgxb;
	output	[1:0]  rx_ctrldetect;
	output	[15:0]  rx_dataout;
	output	[0:0]  rx_freqlocked;
	output	[1:0]  rx_patterndetect;
	output	[0:0]  rx_pll_locked;
	output	[1:0]  rx_syncstatus;
	output	[0:0]  tx_clkout;
	output	[0:0]  tx_dataout;

	parameter		starting_channel_number = 0;


	wire [1:0] sub_wire0;
	wire [1:0] sub_wire1;
	wire [0:0] sub_wire2;
	wire [0:0] sub_wire3;
	wire [0:0] sub_wire4;
	wire [0:0] sub_wire5;
	wire [0:0] sub_wire6;
	wire [0:0] sub_wire7;
	wire [2:0] sub_wire8;
	wire [1:0] sub_wire9;
	wire [0:0] sub_wire10;
	wire [0:0] sub_wire11;
	wire [0:0] sub_wire12;
	wire [15:0] sub_wire13;
	wire [1:0] rx_patterndetect = sub_wire0[1:0];
	wire [1:0] rx_ctrldetect = sub_wire1[1:0];
	wire [0:0] pipedatavalid = sub_wire2[0:0];
	wire [0:0] pipephydonestatus = sub_wire3[0:0];
	wire [0:0] rx_pll_locked = sub_wire4[0:0];
	wire [0:0] rx_freqlocked = sub_wire5[0:0];
	wire [0:0] tx_dataout = sub_wire6[0:0];
	wire [0:0] pipeelecidle = sub_wire7[0:0];
	wire [2:0] pipestatus = sub_wire8[2:0];
	wire [1:0] rx_syncstatus = sub_wire9[1:0];
	wire [0:0] tx_clkout = sub_wire10[0:0];
	wire [0:0] reconfig_fromgxb = sub_wire11[0:0];
	wire [0:0] pll_locked = sub_wire12[0:0];
	wire [15:0] rx_dataout = sub_wire13[15:0];

	alt2gxb	alt2gxb_component (
				.tx_forceelecidle (tx_forceelecidle),
				.pll_inclk (pll_inclk),
				.gxb_powerdown (gxb_powerdown),
				.tx_datain (tx_datain),
				.rx_cruclk (rx_cruclk),
				.cal_blk_clk (cal_blk_clk),
				.powerdn (powerdn),
				.reconfig_clk (reconfig_clk),
				.fixedclk (fixedclk),
				.rx_datain (rx_datain),
				.reconfig_togxb (reconfig_togxb),
				.tx_ctrlenable (tx_ctrlenable),
				.rx_analogreset (rx_analogreset),
				.pipe8b10binvpolarity (pipe8b10binvpolarity),
				.rx_digitalreset (rx_digitalreset),
				.tx_digitalreset (tx_digitalreset),
				.tx_forcedispcompliance (tx_forcedispcompliance),
				.tx_detectrxloop (tx_detectrxloop),
				.rx_patterndetect (sub_wire0),
				.rx_ctrldetect (sub_wire1),
				.pipedatavalid (sub_wire2),
				.pipephydonestatus (sub_wire3),
				.rx_pll_locked (sub_wire4),
				.rx_freqlocked (sub_wire5),
				.tx_dataout (sub_wire6),
				.pipeelecidle (sub_wire7),
				.pipestatus (sub_wire8),
				.rx_syncstatus (sub_wire9),
				.tx_clkout (sub_wire10),
				.reconfig_fromgxb (sub_wire11),
				.pll_locked (sub_wire12),
				.rx_dataout (sub_wire13)
				// synopsys translate_off
				,
				.cal_blk_calibrationstatus (),
				.cal_blk_powerdown (),
				.coreclkout (),
				.debug_rx_phase_comp_fifo_error (),
				.debug_tx_phase_comp_fifo_error (),
				.gxb_enable (),
				.pll_inclk_alt (),
				.pll_locked_alt (),
				.reconfig_fromgxb_oe (),
				.rx_a1a2size (),
				.rx_a1a2sizeout (),
				.rx_a1detect (),
				.rx_a2detect (),
				.rx_bistdone (),
				.rx_bisterr (),
				.rx_bitslip (),
				.rx_byteorderalignstatus (),
				.rx_channelaligned (),
				.rx_clkout (),
				.rx_coreclk (),
				.rx_cruclk_alt (),
				.rx_dataoutfull (),
				.rx_disperr (),
				.rx_enabyteord (),
				.rx_enapatternalign (),
				.rx_errdetect (),
				.rx_invpolarity (),
				.rx_k1detect (),
				.rx_k2detect (),
				.rx_locktodata (),
				.rx_locktorefclk (),
				.rx_phfifooverflow (),
				.rx_phfifordenable (),
				.rx_phfiforeset (),
				.rx_phfifounderflow (),
				.rx_phfifowrdisable (),
				.rx_powerdown (),
				.rx_recovclkout (),
				.rx_revbitorderwa (),
				.rx_revbyteorderwa (),
				.rx_rlv (),
				.rx_rmfifoalmostempty (),
				.rx_rmfifoalmostfull (),
				.rx_rmfifodatadeleted (),
				.rx_rmfifodatainserted (),
				.rx_rmfifoempty (),
				.rx_rmfifofull (),
				.rx_rmfifordena (),
				.rx_rmfiforeset (),
				.rx_rmfifowrena (),
				.rx_runningdisp (),
				.rx_seriallpbken (),
				.rx_signaldetect (),
				.tx_coreclk (),
				.tx_datainfull (),
				.tx_dispval (),
				.tx_forcedisp (),
				.tx_invpolarity (),
				.tx_phfifooverflow (),
				.tx_phfiforeset (),
				.tx_phfifounderflow (),
				.tx_revparallellpbken ()
				// synopsys translate_on
				);
	defparam
		alt2gxb_component.starting_channel_number = starting_channel_number,
		alt2gxb_component.cmu_pll_inclock_period = 10000,
		alt2gxb_component.cmu_pll_loop_filter_resistor_control = 3,
		alt2gxb_component.digitalreset_port_width = 1,
		alt2gxb_component.enable_fast_recovery_pci_mode = "true",
		alt2gxb_component.en_local_clk_div_ctrl = "true",
		alt2gxb_component.equalizer_ctrl_a_setting = 0,
		alt2gxb_component.equalizer_ctrl_b_setting = 0,
		alt2gxb_component.equalizer_ctrl_c_setting = 0,
		alt2gxb_component.equalizer_ctrl_d_setting = 0,
		alt2gxb_component.equalizer_ctrl_v_setting = 0,
		alt2gxb_component.equalizer_dcgain_setting = 1,
		alt2gxb_component.gen_reconfig_pll = "false",
		alt2gxb_component.loopback_mode = "none",
		alt2gxb_component.lpm_type = "alt2gxb",
		alt2gxb_component.number_of_channels = 1,
		alt2gxb_component.operation_mode = "duplex",
		alt2gxb_component.preemphasis_ctrl_1stposttap_setting = 5,
		alt2gxb_component.preemphasis_ctrl_2ndposttap_inv_setting = "false",
		alt2gxb_component.preemphasis_ctrl_2ndposttap_setting = 0,
		alt2gxb_component.preemphasis_ctrl_pretap_inv_setting = "false",
		alt2gxb_component.preemphasis_ctrl_pretap_setting = 0,
		alt2gxb_component.protocol = "pipe",
		alt2gxb_component.receiver_termination = "oct_100_ohms",
		alt2gxb_component.reconfig_dprio_mode = 1,
		alt2gxb_component.reverse_loopback_mode = "rplb",
		alt2gxb_component.rx_8b_10b_compatibility_mode = "true",
		alt2gxb_component.rx_8b_10b_mode = "normal",
		alt2gxb_component.rx_align_pattern = "0101111100",
		alt2gxb_component.rx_align_pattern_length = 10,
		alt2gxb_component.rx_allow_align_polarity_inversion = "false",
		alt2gxb_component.rx_allow_pipe_polarity_inversion = "true",
		alt2gxb_component.rx_bandwidth_mode = 1,
		alt2gxb_component.rx_bitslip_enable = "false",
		alt2gxb_component.rx_byte_ordering_mode = "none",
		alt2gxb_component.rx_channel_bonding = "indv",
		alt2gxb_component.rx_channel_width = 16,
		alt2gxb_component.rx_common_mode = "0.9v",
		alt2gxb_component.rx_cru_inclock_period = 10000,
		alt2gxb_component.rx_cru_pre_divide_by = 1,
		alt2gxb_component.rx_datapath_protocol = "pipe",
		alt2gxb_component.rx_data_rate = 2500,
		alt2gxb_component.rx_data_rate_remainder = 0,
		alt2gxb_component.rx_disable_auto_idle_insertion = "false",
		alt2gxb_component.rx_enable_bit_reversal = "false",
		alt2gxb_component.rx_enable_lock_to_data_sig = "false",
		alt2gxb_component.rx_enable_lock_to_refclk_sig = "false",
		alt2gxb_component.rx_enable_self_test_mode = "false",
		alt2gxb_component.rx_enable_true_complement_match_in_word_align = "false",
		alt2gxb_component.rx_force_signal_detect = "false",
		alt2gxb_component.rx_ppmselect = 8,
		alt2gxb_component.rx_rate_match_back_to_back = "false",
		alt2gxb_component.rx_rate_match_fifo_mode = "normal",
		alt2gxb_component.rx_rate_match_ordered_set_based = "false",
		alt2gxb_component.rx_rate_match_pattern1 = "11010000111010000011",
		alt2gxb_component.rx_rate_match_pattern2 = "00101111000101111100",
		alt2gxb_component.rx_rate_match_pattern_size = 20,
		alt2gxb_component.rx_rate_match_skip_set_based = "false",
		alt2gxb_component.rx_run_length_enable = "false",
		alt2gxb_component.rx_signal_detect_threshold = 1,
		alt2gxb_component.rx_use_align_state_machine = "true",
		alt2gxb_component.rx_use_clkout = "false",
		alt2gxb_component.rx_use_coreclk = "false",
		alt2gxb_component.rx_use_cruclk = "true",
		alt2gxb_component.rx_use_deserializer_double_data_mode = "false",
		alt2gxb_component.rx_use_deskew_fifo = "false",
		alt2gxb_component.rx_use_double_data_mode = "true",
		alt2gxb_component.rx_use_pipe8b10binvpolarity = "true",
		alt2gxb_component.rx_use_rate_match_pattern1_only = "false",
		alt2gxb_component.transmitter_termination = "oct_100_ohms",
		alt2gxb_component.tx_8b_10b_compatibility_mode = "true",
		alt2gxb_component.tx_8b_10b_mode = "normal",
		alt2gxb_component.tx_allow_polarity_inversion = "false",
		alt2gxb_component.tx_analog_power = "1.2v",
		alt2gxb_component.tx_channel_bonding = "indv",
		alt2gxb_component.tx_channel_width = 16,
		alt2gxb_component.tx_common_mode = "0.6v",
		alt2gxb_component.tx_data_rate = 2500,
		alt2gxb_component.tx_data_rate_remainder = 0,
		alt2gxb_component.tx_enable_bit_reversal = "false",
		alt2gxb_component.tx_enable_idle_selection = "false",
		alt2gxb_component.tx_enable_self_test_mode = "false",
		alt2gxb_component.tx_refclk_divide_by = 1,
		alt2gxb_component.tx_transmit_protocol = "pipe",
		alt2gxb_component.tx_use_coreclk = "false",
		alt2gxb_component.tx_use_double_data_mode = "true",
		alt2gxb_component.tx_use_serializer_double_data_mode = "false",
		alt2gxb_component.use_calibration_block = "true",
		alt2gxb_component.vod_ctrl_setting = 4;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ALT_SIMLIB_GEN STRING "0"
// Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
// Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
// Retrieval info: PRIVATE: RX_FORCE_SIGNAL_DETECT STRING "false"
// Retrieval info: PRIVATE: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "1"
// Retrieval info: PRIVATE: VOD_CTRL_SETTING NUMERIC "800"
// Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2500.0000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "62.2"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2500"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "62.2"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "1"
// Retrieval info: PRIVATE: WIZ_EXTERNAL_RX_TERMINATION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_EXTERNAL_TX_TERMINATION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "100"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "100"
// Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2500.0000"
// Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_INPUT_B STRING "100"
// Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "5"
// Retrieval info: PRIVATE: WIZ_PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "PCI Express (PIPE)"
// Retrieval info: PRIVATE: WIZ_RX_TERMINATION NUMERIC "100"
// Retrieval info: PRIVATE: WIZ_RX_VCM STRING "0.85"
// Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "x1"
// Retrieval info: PRIVATE: WIZ_TCL_KEY STRING "STRATIXIIGX_CONFIG_MODE_PIPE_1X"
// Retrieval info: PRIVATE: WIZ_TX_TERMINATION NUMERIC "100"
// Retrieval info: PRIVATE: WIZ_TX_VCM STRING "0.6"
// Retrieval info: PRIVATE: WIZ_VCCHTX STRING "1.2"
// Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
// Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
// Retrieval info: CONSTANT: CMU_PLL_INCLOCK_PERIOD NUMERIC "10000"
// Retrieval info: CONSTANT: CMU_PLL_LOOP_FILTER_RESISTOR_CONTROL NUMERIC "3"
// Retrieval info: CONSTANT: DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: ENABLE_FAST_RECOVERY_PCI_MODE STRING "true"
// Retrieval info: CONSTANT: EN_LOCAL_CLK_DIV_CTRL STRING "true"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_A_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_B_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_C_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_D_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_V_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "1"
// Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
// Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alt2gxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "5"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_INV_SETTING STRING "false"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_INV_SETTING STRING "false"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PROTOCOL STRING "pipe"
// Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "1"
// Retrieval info: CONSTANT: REVERSE_LOOPBACK_MODE STRING "rplb"
// Retrieval info: CONSTANT: RX_8B_10B_COMPATIBILITY_MODE STRING "true"
// Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "normal"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
// Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "true"
// Retrieval info: CONSTANT: RX_BANDWIDTH_MODE NUMERIC "1"
// Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
// Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "none"
// Retrieval info: CONSTANT: RX_CHANNEL_BONDING STRING "indv"
// Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "16"
// Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.9v"
// Retrieval info: CONSTANT: RX_CRU_INCLOCK_PERIOD NUMERIC "10000"
// Retrieval info: CONSTANT: RX_CRU_PRE_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "pipe"
// Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "2500"
// Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: RX_DISABLE_AUTO_IDLE_INSERTION STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_TRUE_COMPLEMENT_MATCH_IN_WORD_ALIGN STRING "false"
// Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "false"
// Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "8"
// Retrieval info: CONSTANT: RX_RATE_MATCH_BACK_TO_BACK STRING "false"
// Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "normal"
// Retrieval info: CONSTANT: RX_RATE_MATCH_ORDERED_SET_BASED STRING "false"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN1 STRING "11010000111010000011"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN2 STRING "00101111000101111100"
// Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN_SIZE NUMERIC "20"
// Retrieval info: CONSTANT: RX_RATE_MATCH_SKIP_SET_BASED STRING "false"
// Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "false"
// Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "1"
// Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "true"
// Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "false"
// Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: RX_USE_CRUCLK STRING "true"
// Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
// Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "true"
// Retrieval info: CONSTANT: RX_USE_PIPE8B10BINVPOLARITY STRING "true"
// Retrieval info: CONSTANT: RX_USE_RATE_MATCH_PATTERN1_ONLY STRING "false"
// Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: TX_8B_10B_COMPATIBILITY_MODE STRING "true"
// Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
// Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "1.2v"
// Retrieval info: CONSTANT: TX_CHANNEL_BONDING STRING "indv"
// Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "16"
// Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.6v"
// Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2500"
// Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: TX_ENABLE_IDLE_SELECTION STRING "false"
// Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: TX_REFCLK_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "pipe"
// Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
// Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
// Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "4"
// Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
// Retrieval info: USED_PORT: fixedclk 0 0 0 0 INPUT NODEFVAL "fixedclk"
// Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
// Retrieval info: USED_PORT: pipe8b10binvpolarity 0 0 1 0 INPUT NODEFVAL "pipe8b10binvpolarity[0..0]"
// Retrieval info: USED_PORT: pipedatavalid 0 0 1 0 OUTPUT NODEFVAL "pipedatavalid[0..0]"
// Retrieval info: USED_PORT: pipeelecidle 0 0 1 0 OUTPUT NODEFVAL "pipeelecidle[0..0]"
// Retrieval info: USED_PORT: pipephydonestatus 0 0 1 0 OUTPUT NODEFVAL "pipephydonestatus[0..0]"
// Retrieval info: USED_PORT: pipestatus 0 0 3 0 OUTPUT NODEFVAL "pipestatus[2..0]"
// Retrieval info: USED_PORT: pll_inclk 0 0 0 0 INPUT NODEFVAL "pll_inclk"
// Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
// Retrieval info: USED_PORT: powerdn 0 0 2 0 INPUT NODEFVAL "powerdn[1..0]"
// Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
// Retrieval info: USED_PORT: reconfig_fromgxb 0 0 1 0 OUTPUT NODEFVAL "reconfig_fromgxb[0..0]"
// Retrieval info: USED_PORT: reconfig_togxb 0 0 3 0 INPUT NODEFVAL "reconfig_togxb[2..0]"
// Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
// Retrieval info: USED_PORT: rx_cruclk 0 0 1 0 INPUT GND "rx_cruclk[0..0]"
// Retrieval info: USED_PORT: rx_ctrldetect 0 0 2 0 OUTPUT NODEFVAL "rx_ctrldetect[1..0]"
// Retrieval info: USED_PORT: rx_datain 0 0 1 0 INPUT NODEFVAL "rx_datain[0..0]"
// Retrieval info: USED_PORT: rx_dataout 0 0 16 0 OUTPUT NODEFVAL "rx_dataout[15..0]"
// Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
// Retrieval info: USED_PORT: rx_freqlocked 0 0 1 0 OUTPUT NODEFVAL "rx_freqlocked[0..0]"
// Retrieval info: USED_PORT: rx_patterndetect 0 0 2 0 OUTPUT NODEFVAL "rx_patterndetect[1..0]"
// Retrieval info: USED_PORT: rx_pll_locked 0 0 1 0 OUTPUT NODEFVAL "rx_pll_locked[0..0]"
// Retrieval info: USED_PORT: rx_syncstatus 0 0 2 0 OUTPUT NODEFVAL "rx_syncstatus[1..0]"
// Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
// Retrieval info: USED_PORT: tx_ctrlenable 0 0 2 0 INPUT NODEFVAL "tx_ctrlenable[1..0]"
// Retrieval info: USED_PORT: tx_datain 0 0 16 0 INPUT NODEFVAL "tx_datain[15..0]"
// Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
// Retrieval info: USED_PORT: tx_detectrxloop 0 0 1 0 INPUT NODEFVAL "tx_detectrxloop[0..0]"
// Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
// Retrieval info: USED_PORT: tx_forcedispcompliance 0 0 1 0 INPUT NODEFVAL "tx_forcedispcompliance[0..0]"
// Retrieval info: USED_PORT: tx_forceelecidle 0 0 1 0 INPUT NODEFVAL "tx_forceelecidle[0..0]"
// Retrieval info: CONNECT: @fixedclk 0 0 0 0 fixedclk 0 0 0 0
// Retrieval info: CONNECT: @tx_detectrxloop 0 0 1 0 tx_detectrxloop 0 0 1 0
// Retrieval info: CONNECT: @tx_forcedispcompliance 0 0 1 0 tx_forcedispcompliance 0 0 1 0
// Retrieval info: CONNECT: rx_patterndetect 0 0 2 0 @rx_patterndetect 0 0 2 0
// Retrieval info: CONNECT: pipedatavalid 0 0 1 0 @pipedatavalid 0 0 1 0
// Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
// Retrieval info: CONNECT: @powerdn 0 0 2 0 powerdn 0 0 2 0
// Retrieval info: CONNECT: pipeelecidle 0 0 1 0 @pipeelecidle 0 0 1 0
// Retrieval info: CONNECT: rx_ctrldetect 0 0 2 0 @rx_ctrldetect 0 0 2 0
// Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
// Retrieval info: CONNECT: rx_dataout 0 0 16 0 @rx_dataout 0 0 16 0
// Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
// Retrieval info: CONNECT: pipestatus 0 0 3 0 @pipestatus 0 0 3 0
// Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: rx_pll_locked 0 0 1 0 @rx_pll_locked 0 0 1 0
// Retrieval info: CONNECT: rx_syncstatus 0 0 2 0 @rx_syncstatus 0 0 2 0
// Retrieval info: CONNECT: @pipe8b10binvpolarity 0 0 1 0 pipe8b10binvpolarity 0 0 1 0
// Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
// Retrieval info: CONNECT: @reconfig_togxb 0 0 3 0 reconfig_togxb 0 0 3 0
// Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
// Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
// Retrieval info: CONNECT: @rx_cruclk 0 0 1 0 rx_cruclk 0 0 1 0
// Retrieval info: CONNECT: @pll_inclk 0 0 0 0 pll_inclk 0 0 0 0
// Retrieval info: CONNECT: @tx_ctrlenable 0 0 2 0 tx_ctrlenable 0 0 2 0
// Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
// Retrieval info: CONNECT: @tx_datain 0 0 16 0 tx_datain 0 0 16 0
// Retrieval info: CONNECT: reconfig_fromgxb 0 0 1 0 @reconfig_fromgxb 0 0 1 0
// Retrieval info: CONNECT: rx_freqlocked 0 0 1 0 @rx_freqlocked 0 0 1 0
// Retrieval info: CONNECT: @rx_datain 0 0 1 0 rx_datain 0 0 1 0
// Retrieval info: CONNECT: pipephydonestatus 0 0 1 0 @pipephydonestatus 0 0 1 0
// Retrieval info: CONNECT: @tx_forceelecidle 0 0 1 0 tx_forceelecidle 0 0 1 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_serdes_2sgx_x1d_10000_bb.v FALSE FALSE
