-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt2gxb_reconfig 

-- ============================================================
-- File Name: altpcie_reconfig_4sgx.vhd
-- Megafunction Name(s):
-- 			alt2gxb_reconfig
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Internal Build 134 03/09/2011 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt2gxb_reconfig BASE_PORT_WIDTH=1 CBX_AUTO_BLACKBOX="ALL" CHANNEL_ADDRESS_WIDTH=3 DEVICE_FAMILY="Stratix IV" ENABLE_BUF_CAL="TRUE" ENABLE_CHL_ADDR_FOR_ANALOG_CTRL="TRUE" NUMBER_OF_CHANNELS=8 NUMBER_OF_RECONFIG_PORTS=2 READ_BASE_PORT_WIDTH=1 RECONFIG_FROMGXB_WIDTH=34 RECONFIG_TOGXB_WIDTH=4 RX_EQDCGAIN_PORT_WIDTH=3 TX_PREEMP_PORT_WIDTH=5 busy data_valid logical_channel_address offset_cancellation_reset read reconfig_clk reconfig_fromgxb reconfig_mode_sel reconfig_togxb rx_eqctrl rx_eqctrl_out rx_eqdcgain rx_eqdcgain_out tx_preemp_0t tx_preemp_0t_out tx_preemp_1t tx_preemp_1t_out tx_preemp_2t tx_preemp_2t_out tx_vodctrl tx_vodctrl_out write_all
--VERSION_BEGIN 11.0 cbx_alt2gxb_reconfig 2011:03:09:22:37:51:SJ cbx_alt_cal 2011:03:09:22:37:51:SJ cbx_alt_dprio 2011:03:09:22:37:51:SJ cbx_altsyncram 2011:03:09:22:37:54:SJ cbx_cycloneii 2011:03:09:22:37:55:SJ cbx_lpm_add_sub 2011:03:09:22:37:56:SJ cbx_lpm_compare 2011:03:09:22:37:56:SJ cbx_lpm_counter 2011:03:09:22:37:56:SJ cbx_lpm_decode 2011:03:09:22:37:56:SJ cbx_lpm_mux 2011:03:09:22:37:56:SJ cbx_lpm_shiftreg 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ cbx_stratix 2011:03:09:22:37:58:SJ cbx_stratixii 2011:03:09:22:37:58:SJ cbx_stratixiii 2011:03:09:22:37:58:SJ cbx_stratixv 2011:03:09:22:37:58:SJ cbx_util_mgl 2011:03:09:22:37:57:SJ  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Stratix IV" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset wren wren_data
--VERSION_BEGIN 11.0 cbx_alt_dprio 2011:03:09:22:37:51:SJ cbx_cycloneii 2011:03:09:22:37:55:SJ cbx_lpm_add_sub 2011:03:09:22:37:56:SJ cbx_lpm_compare 2011:03:09:22:37:56:SJ cbx_lpm_counter 2011:03:09:22:37:56:SJ cbx_lpm_decode 2011:03:09:22:37:56:SJ cbx_lpm_shiftreg 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ cbx_stratix 2011:03:09:22:37:58:SJ cbx_stratixii 2011:03:09:22:37:58:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_4sgx_alt_dprio_2vj IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END altpcie_reconfig_4sgx_alt_dprio_2vj;

 ARCHITECTURE RTL OF altpcie_reconfig_4sgx_alt_dprio_2vj IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1191w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1195w1201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1195w1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1187w1188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1187w1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1187w1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1195w1196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range1061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb948w1125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb948w1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_0787w788w789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_0806w807w808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_0822w823w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren776w799w812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren776w799w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state947w951w952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state1127w1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state1062w1063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_0787w788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_0806w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_0822w823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren776w799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren776w777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren776w794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1183w1184w1185w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state947w951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state1127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state1062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_0787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_0806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_0822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden1183w1184w1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden774w775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1183w1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_1790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_1809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_1825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_0787w788w789w(0) <= wire_dprio_w_lg_w_lg_s0_to_0787w788w(0) AND wire_state_mc_reg_w_q_range785w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_0806w807w808w(0) <= wire_dprio_w_lg_w_lg_s1_to_0806w807w(0) AND wire_state_mc_reg_w_q_range804w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_0822w823w824w(0) <= wire_dprio_w_lg_w_lg_s2_to_0822w823w(0) AND wire_state_mc_reg_w_q_range820w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren776w799w812w(0) <= wire_dprio_w_lg_w_lg_wren776w799w(0) AND wire_dprio_w_lg_rdinc811w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren776w799w800w(0) <= wire_dprio_w_lg_w_lg_wren776w799w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state947w951w952w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state947w951w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state1127w1128w(0) <= wire_dprio_w_lg_rd_data_output_state1127w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state1062w1063w(0) <= wire_dprio_w_lg_wr_data_state1062w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_0787w788w(0) <= wire_dprio_w_lg_s0_to_0787w(0) AND wire_dprio_w_lg_s0_to_1786w(0);
	wire_dprio_w_lg_w_lg_s1_to_0806w807w(0) <= wire_dprio_w_lg_s1_to_0806w(0) AND wire_dprio_w_lg_s1_to_1805w(0);
	wire_dprio_w_lg_w_lg_s2_to_0822w823w(0) <= wire_dprio_w_lg_s2_to_0822w(0) AND wire_dprio_w_lg_s2_to_1821w(0);
	wire_dprio_w_lg_w_lg_wren776w799w(0) <= wire_dprio_w_lg_wren776w(0) AND wire_dprio_w_lg_wren_data798w(0);
	wire_dprio_w_lg_w_lg_wren776w777w(0) <= wire_dprio_w_lg_wren776w(0) AND wire_dprio_w_lg_w_lg_rden774w775w(0);
	wire_dprio_w_lg_w_lg_wren776w794w(0) <= wire_dprio_w_lg_wren776w(0) AND wire_dprio_w_lg_rdinc793w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1183w1184w1185w1186w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden1183w1184w1185w(0) AND wire_dprio_w_lg_startup_done1181w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state947w951w(0) <= wire_dprio_w_lg_wr_addr_state947w(0) AND wire_addr_shift_reg_w_q_range950w(0);
	wire_dprio_w_lg_idle_state813w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren776w799w812w(0);
	wire_dprio_w_lg_idle_state795w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren776w794w(0);
	wire_dprio_w_lg_idle_state802w(0) <= idle_state AND wire_dprio_w_lg_wren801w(0);
	wire_dprio_w_lg_idle_state779w(0) <= idle_state AND wire_dprio_w_lg_wren778w(0);
	wire_dprio_w_lg_idle_state816w(0) <= idle_state AND wire_dprio_w_lg_wren815w(0);
	wire_dprio_w_lg_rd_data_output_state1127w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range1126w(0);
	wire_dprio_w_lg_wr_data_state1062w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range1061w(0);
	wire_dprio_w_lg_s0_to_0787w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_1786w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_0806w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_1805w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_0822w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_1821w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done1181w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle1182w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren776w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data798w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden1183w1184w1185w(0) <= wire_dprio_w_lg_w_lg_rden1183w1184w(0) OR wire_dprio_w_lg_startup_idle1182w(0);
	wire_dprio_w_lg_w_lg_rden774w775w(0) <= wire_dprio_w_lg_rden774w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden1183w1184w(0) <= wire_dprio_w_lg_rden1183w(0) OR rdinc;
	wire_dprio_w_lg_rden774w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden1183w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc811w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc793w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_1790w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_0787w788w789w(0);
	wire_dprio_w_lg_s1_to_1809w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_0806w807w808w(0);
	wire_dprio_w_lg_s2_to_1825w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_0822w823w824w(0);
	wire_dprio_w_lg_wr_addr_state947w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren801w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren776w799w800w(0);
	wire_dprio_w_lg_wren778w(0) <= wren OR wire_dprio_w_lg_w_lg_wren776w777w(0);
	wire_dprio_w_lg_wren815w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range1195w1204w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range1187w1192w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state779w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state802w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state795w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state816w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state813w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range1195w1201w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range1187w1188w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range950w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range1126w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range1195w1196w & wire_startup_cntr_w_lg_w_q_range1187w1192w & wire_startup_cntr_w_lg_w_q_range1187w1188w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1183w1184w1185w1186w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range1191w1194w(0) <= wire_startup_cntr_w_q_range1191w(0) AND wire_startup_cntr_w_q_range1187w(0);
	wire_startup_cntr_w_lg_w_q_range1195w1201w(0) <= wire_startup_cntr_w_q_range1195w(0) AND wire_startup_cntr_w_lg_w_q_range1187w1188w(0);
	wire_startup_cntr_w_lg_w_q_range1195w1204w(0) <= wire_startup_cntr_w_q_range1195w(0) AND wire_startup_cntr_w_lg_w_q_range1187w1203w(0);
	wire_startup_cntr_w_lg_w_q_range1187w1188w(0) <= NOT wire_startup_cntr_w_q_range1187w(0);
	wire_startup_cntr_w_lg_w_q_range1187w1203w(0) <= wire_startup_cntr_w_q_range1187w(0) OR wire_startup_cntr_w_q_range1191w(0);
	wire_startup_cntr_w_lg_w_q_range1187w1192w(0) <= wire_startup_cntr_w_q_range1187w(0) XOR wire_startup_cntr_w_q_range1191w(0);
	wire_startup_cntr_w_lg_w_q_range1195w1196w(0) <= wire_startup_cntr_w_q_range1195w(0) XOR wire_startup_cntr_w_lg_w_q_range1191w1194w(0);
	wire_startup_cntr_w_q_range1187w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range1191w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range1195w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_1825w & wire_dprio_w_lg_s1_to_1809w & wire_dprio_w_lg_s0_to_1790w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range785w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range804w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range820w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range1061w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb948w1125w(0) <= wire_pre_amble_cmpr_w_lg_agb948w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb948w1060w(0) <= wire_pre_amble_cmpr_w_lg_agb948w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb948w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state770w(0);
	wire_dprio_w_lg_write_state770w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state947w951w952w(0) OR (wire_pre_amble_cmpr_w_lg_agb948w(0) AND wire_dprio_w_lg_wr_addr_state947w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state1062w1063w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb948w1060w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state1127w1128w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb948w1125w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --altpcie_reconfig_4sgx_alt_dprio_2vj


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=8 LPM_WIDTH=1 LPM_WIDTHS=3 data result sel
--VERSION_BEGIN 11.0 cbx_lpm_mux 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ  VERSION_END

--synthesis_resources = lut 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_4sgx_mux_c6a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altpcie_reconfig_4sgx_mux_c6a;

 ARCHITECTURE RTL OF altpcie_reconfig_4sgx_mux_c6a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l2_w0_n1_mux_dataout & wire_l2_w0_n0_mux_dataout & wire_l1_w0_n3_mux_dataout & wire_l1_w0_n2_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & data);
	result <= result_wire_ext;
	result_wire_ext(0) <= ( wire_l3_w0_n0_mux_dataout);
	sel_wire <= ( sel(2) & "000" & sel(1) & "000" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(1) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(3) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w0_n2_mux_dataout <= data_wire(5) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w0_n3_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(6);
	wire_l2_w0_n0_mux_dataout <= data_wire(9) WHEN sel_wire(4) = '1'  ELSE data_wire(8);
	wire_l2_w0_n1_mux_dataout <= data_wire(11) WHEN sel_wire(4) = '1'  ELSE data_wire(10);
	wire_l3_w0_n0_mux_dataout <= data_wire(13) WHEN sel_wire(8) = '1'  ELSE data_wire(12);

 END RTL; --altpcie_reconfig_4sgx_mux_c6a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=2 LPM_WIDTH=1 LPM_WIDTHS=1 data result sel
--VERSION_BEGIN 11.0 cbx_lpm_mux 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ  VERSION_END

--synthesis_resources = lut 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_4sgx_mux_46a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END altpcie_reconfig_4sgx_mux_46a;

 ARCHITECTURE RTL OF altpcie_reconfig_4sgx_mux_46a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	data_wire <= ( data);
	result <= result_wire_ext;
	result_wire_ext(0) <= ( wire_l1_w0_n0_mux_dataout);
	sel_wire(0) <= ( sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(1) WHEN sel_wire(0) = '1'  ELSE data_wire(0);

 END RTL; --altpcie_reconfig_4sgx_mux_46a

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = alt_cal 1 lpm_add_sub 4 lpm_compare 7 lpm_counter 4 lpm_decode 3 lut 5 reg 149 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 logical_channel_address	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 offset_cancellation_reset	:	IN  STD_LOGIC := '0';
		 read	:	IN  STD_LOGIC := '0';
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 reconfig_mode_sel	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_eqctrl	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 rx_eqctrl_out	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_eqdcgain	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 rx_eqdcgain_out	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 tx_preemp_0t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_0t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_preemp_1t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_1t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_preemp_2t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_2t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_vodctrl	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 tx_vodctrl_out	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 write_all	:	IN  STD_LOGIC := '0'
	 ); 
 END altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1;

 ARCHITECTURE RTL OF altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0";

	 SIGNAL  wire_calibration_w_lg_w_lg_busy171w175w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy171w172w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy171w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy171w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy171w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy176w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy173w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range704w705w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range704w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range704w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range497w706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range497w716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range688w689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_busy199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range684w687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range707w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range704w705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_dataout_range704w705w717w718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range704w713w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range704w708w709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_dataout_range692w693w694w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range692w693w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range692w693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy176w177w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy173w174w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy179w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren_data	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy185w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range410w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range730w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range742w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_q_range136w137w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range140w141w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range136w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range136w137w138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range140w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 data_valid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF data_valid_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_data_valid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 dprio_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 reconf_mode_sel_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconf_mode_sel_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rx_eqctrl_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 rx_eqctrl_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rx_eqctrl_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rx_eqctrl_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_rx_equalizer_dcgain_reg_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 rx_equalizer_dcgain_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rx_equalizer_dcgain_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rx_equalizer_dcgain_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := "00"
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_lg_q31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_lg_q29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tx_preemp_0t_inv_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemp_0t_inv_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemp_0t_inv_reg_ena	:	STD_LOGIC_VECTOR(0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_0t_inv_reg_w_lg_w_q_range752w753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_0t_inv_reg_w_q_range752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tx_preemp_2t_inv_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemp_2t_inv_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemp_2t_inv_reg_ena	:	STD_LOGIC_VECTOR(0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_2t_inv_reg_w_lg_w_q_range762w763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_2t_inv_reg_w_q_range762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_1stposttap_reg_d	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_1stposttap_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_1stposttap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_1stposttap_reg_ena	:	STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_2ndposttap_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_2ndposttap_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_2ndposttap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_2ndposttap_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_pretap_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_pretap_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_pretap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_pretap_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_tx_vodctrl_reg_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 tx_vodctrl_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_vodctrl_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_vodctrl_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 wr_addr_inc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_addr_inc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_rd_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_rd_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wr_rd_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_wr_rd_pulse_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wren_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wren_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wren_data_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_wren_data_reg_w_lg_w_lg_q337w338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub1_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub10_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_add_sub10_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub10_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub11_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_add_sub11_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub11_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub2_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr6_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr6_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr7_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr7_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr8_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr8_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr9_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr9_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_addr_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_write_done256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_idle_state258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range307w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range305w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range305w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range311w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_addr_inc285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_data	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_read_done286w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state295w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range543w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range541w564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range541w544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range547w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range547w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_data	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_write_done523w524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state531w532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_chl_addr_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_aeq_ch_done_mux_result	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprioout_mux_result	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprioout_mux_sel	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy190w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w456w457w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w459w473w474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_header_proc225w226w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_s2_to_058w59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_s2_to_058w70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w463w464w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain348w349w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1246w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_gt_0_577w609w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_done519w520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range453w461w462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range453w484w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w456w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w482w483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w459w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w459w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w459w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range627w646w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w486w487w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy89w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy89w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy89w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy89w90w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_header_proc225w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_global_clk_div9w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig17w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_3313w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s2_to_058w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s2_to_058w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_reconfig_mode_sel_range81w82w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w463w464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range627w632w633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w125w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w365w366w367w368w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_tier_1350w351w352w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_68_6B355w356w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range122w123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range107w108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range119w120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range103w104w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy91w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain348w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_64_67357w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f354w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f_inv353w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_preemp1t360w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_vodctrl362w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_3312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_59102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_61117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address192w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state681w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state701w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state724w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state737w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state731w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state743w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_64_67_data_valid698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_68_6B_data_valid678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_7c_7f_data_valid739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_7c_7f_inv_data_valid316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_preemp_1t_data_valid734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_vodctrl_data_valid721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_0_617w673w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_10_658w670w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_3_639w672w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_6_649w671w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_0_577w605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_0_577w609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_address193w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_all25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state680w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state700w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state736w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state723w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state729w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state741w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_7c_7f_inv_data_valid551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_done519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range451w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range451w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range453w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range453w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range455w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range455w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range455w459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range433w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range374w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range374w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range372w384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range372w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range455w486w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range372w373w381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range624w625w626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range627w654w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bonded_skip237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_header_proc225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_global_clk_div9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr0239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_diff_mif196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_global_clk_div_mode235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_protected_bit236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_3313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rd_pulse143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_done212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_reconf_addr224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rx_reconfig315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s1_to_068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s1_to_169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s2_to_058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tx_reconfig294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_10_595w602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_3_583w604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_6_589w603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_all_int47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_done229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range76w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range81w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range458w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range451w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range453w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range455w463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_preemp_0t_range2w509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_preemp_2t_range4w513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range371w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range623w630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range624w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w489w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_3313w14w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w125w126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy91w92w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy130w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_vodctrl362w363w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state727w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state681w682w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state701w702w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state724w725w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state737w738w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state731w732w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state743w744w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_64_67_data_valid698w699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_68_6B_data_valid678w679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_7c_7f_data_valid739w740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_preemp_1t_data_valid734w735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_vodctrl_data_valid721w722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range451w467w468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range451w477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range372w384w385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range372w376w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig17w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1222w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1222w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w489w490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w110w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl362w363w364w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range451w467w468w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w489w490w491w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w365w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w489w490w491w492w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w365w366w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w470w471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w365w366w367w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w219w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_adce39w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_address95w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s0_to_262w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s0_to_273w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_preemp1t_data_valid358w359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqdcgain_range429w437w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv572w_range627w662w663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_68_6B355w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_adce39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_preemp1t_data_valid358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_vodctrl_data_valid361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range122w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range107w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range119w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range103w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range81w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range429w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range429w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range458w476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range453w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range455w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range372w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range624w625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv572w_range627w654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a2gr_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_rden :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren_data :	STD_LOGIC;
	 SIGNAL  adce_busy_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  aeq_ch_done :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bonded_skip :	STD_LOGIC;
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_channel_address_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  cal_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  channel_address_out :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  dfe_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  diff_mif_wr_rd_busy :	STD_LOGIC;
	 SIGNAL  dprio_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_64_67 :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_68_6B :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f_inv :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_preemp1t :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_vodctrl :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_pulse :	STD_LOGIC;
	 SIGNAL  en_read_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  en_write_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  header_proc :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  internal_write_pulse :	STD_LOGIC;
	 SIGNAL  is_adce :	STD_LOGIC;
	 SIGNAL  is_adce_all_control :	STD_LOGIC;
	 SIGNAL  is_adce_continuous_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_one_time_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_standby_single_control :	STD_LOGIC;
	 SIGNAL  is_analog_control :	STD_LOGIC;
	 SIGNAL  is_bonded_global_clk_div :	STD_LOGIC;
	 SIGNAL  is_bonded_reconfig :	STD_LOGIC;
	 SIGNAL  is_central_pcs :	STD_LOGIC;
	 SIGNAL  is_cruclk_addr0 :	STD_LOGIC;
	 SIGNAL  is_diff_mif :	STD_LOGIC;
	 SIGNAL  is_do_dfe :	STD_LOGIC;
	 SIGNAL  is_do_eyemon :	STD_LOGIC;
	 SIGNAL  is_global_clk_div_mode :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_d :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_out :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  is_pll_address :	STD_LOGIC;
	 SIGNAL  is_protected_bit :	STD_LOGIC;
	 SIGNAL  is_rcxpat_chnl_en_ch :	STD_LOGIC;
	 SIGNAL  is_table_33 :	STD_LOGIC;
	 SIGNAL  is_table_59 :	STD_LOGIC;
	 SIGNAL  is_table_61 :	STD_LOGIC;
	 SIGNAL  is_tier_1 :	STD_LOGIC;
	 SIGNAL  is_tier_2 :	STD_LOGIC;
	 SIGNAL  is_tx_local_div_ctrl :	STD_LOGIC;
	 SIGNAL  legal_rd_mode_type :	STD_LOGIC;
	 SIGNAL  legal_wr_mode_type :	STD_LOGIC;
	 SIGNAL  local_ch_dec :	STD_LOGIC;
	 SIGNAL  logical_pll_sel_num :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  mif_reconfig_done :	STD_LOGIC;
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  quad_address_out :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rd_pulse :	STD_LOGIC;
	 SIGNAL  read_addr_inc :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_done :	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  read_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_7c_7f_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_7c_7f_inv_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_done :	STD_LOGIC;
	 SIGNAL  read_word_preemp_1t_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  reconfig_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 SIGNAL  reset_addr_done :	STD_LOGIC;
	 SIGNAL  reset_reconf_addr :	STD_LOGIC;
	 SIGNAL  reset_system :	STD_LOGIC;
	 SIGNAL  rx_reconfig :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s0_to_2 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  start	:	STD_LOGIC;
	 SIGNAL  state_mc_reg_in :	STD_LOGIC_VECTOR (1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  transceiver_init	:	STD_LOGIC;
	 SIGNAL  tx_preemp_0t_out_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_0t_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_2t_out_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_2t_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_reconfig :	STD_LOGIC;
	 SIGNAL  w334w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  w_eq_0_617w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_10_658w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_3_639w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_6_649w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_gt_0_577w :	STD_LOGIC;
	 SIGNAL  w_gt_0_only601w :	STD_LOGIC;
	 SIGNAL  w_gt_10_595w :	STD_LOGIC;
	 SIGNAL  w_gt_10_only615w :	STD_LOGIC;
	 SIGNAL  w_gt_3_583w :	STD_LOGIC;
	 SIGNAL  w_gt_3_only608w :	STD_LOGIC;
	 SIGNAL  w_gt_6_589w :	STD_LOGIC;
	 SIGNAL  w_gt_6_only612w :	STD_LOGIC;
	 SIGNAL  w_rx_eqa571w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqb570w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqc569w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqctrl_out567w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_rx_eqd568w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqdcgain_out683w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqv572w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_tx_vodctrl_out703w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wr_pulse :	STD_LOGIC;
	 SIGNAL  write_addr_inc :	STD_LOGIC;
	 SIGNAL  write_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_all_int :	STD_LOGIC;
	 SIGNAL  write_done :	STD_LOGIC;
	 SIGNAL  write_happened :	STD_LOGIC;
	 SIGNAL  write_skip :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 SIGNAL  write_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_inv_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_done :	STD_LOGIC;
	 SIGNAL  write_word_preemp1t_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1ta_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1tb_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrla_data_valid :	STD_LOGIC;
	 SIGNAL  wire_w_cal_channel_address_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_channel_address_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_0t_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_0t_wire_range507w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_2t_range4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_2t_wire_range511w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv572w_range623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv572w_range624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv572w_range627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_cal
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "alt_cal"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS*4-1 DOWNTO 0) := (OTHERS => '0');
		transceiver_init	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  altpcie_reconfig_4sgx_alt_dprio_2vj
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altpcie_reconfig_4sgx_mux_c6a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altpcie_reconfig_4sgx_mux_46a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w(0) <= wire_w_lg_w_lg_w_lg_s2_to_058w59w60w(0) AND wire_state_mc_reg_w_q_range55w(0);
	wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w(0) <= wire_w_lg_w_lg_w_lg_s2_to_058w70w71w(0) AND wire_state_mc_reg_w_q_range67w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w456w457w480w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range455w456w457w(0) AND wire_w_rx_eqctrl_range458w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w459w473w474w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range455w459w473w(0) AND wire_w_lg_w_rx_eqctrl_range458w466w(0);
	wire_w489w(0) <= wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w486w487w488w(0) AND wire_w_rx_eqctrl_range458w(0);
	wire_w_lg_w_lg_w_lg_header_proc225w226w227w(0) <= wire_w_lg_w_lg_header_proc225w226w(0) AND wire_w_lg_w_lg_is_tier_1222w223w(0);
	wire_w_lg_w_lg_w_lg_s2_to_058w59w60w(0) <= wire_w_lg_w_lg_s2_to_058w59w(0) AND wire_w_lg_s0_to_056w(0);
	wire_w_lg_w_lg_w_lg_s2_to_058w70w71w(0) <= wire_w_lg_w_lg_s2_to_058w70w(0) AND wire_w_lg_s1_to_068w(0);
	wire_w86w(0) <= wire_w_lg_w_lg_w_reconfig_mode_sel_range81w82w85w(0) AND wire_w_lg_w_reconfig_mode_sel_range76w77w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w463w464w465w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range455w463w464w(0) AND wire_w_rx_eqctrl_range451w(0);
	wire_w634w(0) <= wire_w_lg_w_lg_w_w_rx_eqv572w_range627w632w633w(0) AND wire_w_lg_w_w_rx_eqv572w_range623w630w(0);
	loop1 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain348w349w(i) <= wire_w_lg_dprio_datain348w(i) AND write_state;
	END GENERATE loop1;
	wire_w_lg_w_lg_is_tier_1246w248w(0) <= wire_w_lg_is_tier_1246w(0) AND wire_w_lg_w219w220w(0);
	wire_w_lg_w_lg_w_gt_0_577w609w613w(0) <= wire_w_lg_w_gt_0_577w609w(0) AND w_gt_6_589w;
	wire_w_lg_w_lg_write_word_done519w520w(0) <= wire_w_lg_write_word_done519w(0) AND write_happened;
	wire_w_lg_w_lg_w_rx_eqctrl_range453w461w462w(0) <= wire_w_lg_w_rx_eqctrl_range453w461w(0) AND wire_w_rx_eqctrl_range458w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range453w484w485w(0) <= wire_w_lg_w_rx_eqctrl_range453w484w(0) AND wire_w_lg_w_rx_eqctrl_range458w466w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w456w457w(0) <= wire_w_lg_w_rx_eqctrl_range455w456w(0) AND wire_w_lg_w_rx_eqctrl_range451w452w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w482w483w(0) <= wire_w_lg_w_rx_eqctrl_range455w482w(0) AND wire_w_lg_w_rx_eqctrl_range458w466w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w459w481w(0) <= wire_w_lg_w_rx_eqctrl_range455w459w(0) AND wire_w_lg_w_rx_eqctrl_range458w466w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w459w473w(0) <= wire_w_lg_w_rx_eqctrl_range455w459w(0) AND wire_w_lg_w_rx_eqctrl_range451w452w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w459w460w(0) <= wire_w_lg_w_rx_eqctrl_range455w459w(0) AND wire_w_rx_eqctrl_range458w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range627w646w647w(0) <= wire_w_lg_w_w_rx_eqv572w_range627w646w(0) AND wire_w_lg_w_w_rx_eqv572w_range623w630w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w(0) <= wire_w_lg_w_w_rx_eqv572w_range627w635w(0) AND wire_w_w_rx_eqv572w_range623w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w486w487w488w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range455w486w487w(0) AND wire_w_rx_eqctrl_range451w(0);
	wire_w_lg_w_lg_cal_busy89w128w(0) <= wire_w_lg_cal_busy89w(0) AND wire_w_lg_w_lg_w125w126w127w(0);
	wire_w_lg_w_lg_cal_busy89w112w(0) <= wire_w_lg_cal_busy89w(0) AND wire_w_lg_w110w111w(0);
	wire_w_lg_w_lg_cal_busy89w97w(0) <= wire_w_lg_cal_busy89w(0) AND wire_w_lg_w_lg_is_pll_address95w96w(0);
	loop2 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy89w90w(i) <= wire_w_lg_cal_busy89w(0) AND quad_address(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_header_proc225w226w(0) <= wire_w_lg_header_proc225w(0) AND wire_w_lg_reset_reconf_addr224w(0);
	wire_w_lg_w_lg_is_bonded_global_clk_div9w10w(0) <= wire_w_lg_is_bonded_global_clk_div9w(0) AND busy_state;
	wire_w_lg_w_lg_is_bonded_reconfig17w18w(0) <= wire_w_lg_is_bonded_reconfig17w(0) AND busy_state;
	wire_w_lg_w_lg_is_table_3313w14w(0) <= wire_w_lg_is_table_3313w(0) AND busy_state;
	wire_w_lg_w_lg_s2_to_058w59w(0) <= wire_w_lg_s2_to_058w(0) AND wire_w_lg_s0_to_157w(0);
	wire_w_lg_w_lg_s2_to_058w70w(0) <= wire_w_lg_s2_to_058w(0) AND wire_w_lg_s1_to_169w(0);
	wire_w_lg_w_lg_w_reconfig_mode_sel_range81w82w85w(0) <= wire_w_lg_w_reconfig_mode_sel_range81w82w(0) AND wire_w_reconfig_mode_sel_range78w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w463w464w(0) <= wire_w_lg_w_rx_eqctrl_range455w463w(0) AND wire_w_lg_w_rx_eqctrl_range453w454w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w656w(0) <= wire_w_lg_w_w_rx_eqv572w_range624w631w(0) AND wire_w_lg_w_lg_w_w_rx_eqv572w_range627w654w655w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w667w(0) <= wire_w_lg_w_w_rx_eqv572w_range624w631w(0) AND wire_w_lg_w_w_rx_eqv572w_range623w630w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range627w632w633w(0) <= wire_w_lg_w_w_rx_eqv572w_range627w632w(0) AND wire_w_lg_w_w_rx_eqv572w_range624w631w(0);
	wire_w_lg_w125w126w(0) <= wire_w125w(0) AND wire_w_lg_is_central_pcs118w(0);
	loop3 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_w365w366w367w368w(i) <= wire_w_lg_w_lg_w365w366w367w(i) AND is_analog_control;
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_is_tier_1350w351w352w(i) <= wire_w_lg_w_lg_is_tier_1350w351w(0) AND reconfig_datain(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_68_6B355w356w(i) <= wire_w_lg_dprio_datain_68_6B355w(i) AND write_word_68_6B_data_valid;
	END GENERATE loop5;
	wire_w_lg_w_lg_w_channel_address_range122w123w124w(0) <= wire_w_lg_w_channel_address_range122w123w(0) AND wire_w_lg_is_pll_address106w(0);
	wire_w_lg_w_lg_w_channel_address_range107w108w109w(0) <= wire_w_lg_w_channel_address_range107w108w(0) AND wire_w_lg_is_pll_address106w(0);
	wire_w_lg_w_lg_w_logical_pll_sel_num_range119w120w121w(0) <= wire_w_lg_w_logical_pll_sel_num_range119w120w(0) AND is_pll_address;
	wire_w_lg_w_lg_w_logical_pll_sel_num_range103w104w105w(0) <= wire_w_lg_w_logical_pll_sel_num_range103w104w(0) AND is_pll_address;
	loop6 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_cal_busy91w(i) <= cal_busy AND cal_quad_address(i);
	END GENERATE loop6;
	wire_w_lg_cal_busy130w(0) <= cal_busy AND wire_w_cal_channel_address_range129w(0);
	wire_w_lg_cal_busy114w(0) <= cal_busy AND wire_w_cal_channel_address_range113w(0);
	wire_w_lg_cal_busy99w(0) <= cal_busy AND wire_w_cal_channel_address_range98w(0);
	wire_w_lg_cal_busy190w(0) <= cal_busy AND wire_w_cal_quad_address_range189w(0);
	loop7 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain348w(i) <= dprio_datain(i) AND wire_w_lg_header_proc225w(0);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_64_67357w(i) <= dprio_datain_64_67(i) AND write_word_64_67_data_valid;
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f354w(i) <= dprio_datain_7c_7f(i) AND write_word_7c_7f_data_valid;
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f_inv353w(i) <= dprio_datain_7c_7f_inv(i) AND write_word_7c_7f_inv_data_valid;
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_preemp1t360w(i) <= dprio_datain_preemp1t(i) AND wire_w_lg_w_lg_write_word_preemp1t_data_valid358w359w(0);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_vodctrl362w(i) <= dprio_datain_vodctrl(i) AND wire_w_lg_write_word_vodctrl_data_valid361w(0);
	END GENERATE loop12;
	wire_w_lg_dprio_pulse322w(0) <= dprio_pulse AND wire_read_addr_cntr_w_lg_w_q_range305w321w(0);
	wire_w_lg_dprio_pulse329w(0) <= dprio_pulse AND wire_read_addr_cntr_w_q_range305w(0);
	wire_w_lg_idle_state50w(0) <= idle_state AND wire_w_lg_read49w(0);
	wire_w_lg_idle_state41w(0) <= idle_state AND wire_w_lg_w_lg_is_adce39w40w(0);
	wire_w_lg_is_bonded_reconfig23w(0) <= is_bonded_reconfig AND wire_w_lg_is_bonded_global_clk_div9w(0);
	wire_w_lg_is_bonded_reconfig16w(0) <= is_bonded_reconfig AND wire_w_lg_w_lg_w_lg_is_table_3313w14w15w(0);
	wire_w_lg_is_table_3312w(0) <= is_table_33 AND wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w(0);
	wire_w_lg_is_table_59102w(0) <= is_table_59 AND is_bonded_reconfig;
	wire_w_lg_is_table_61117w(0) <= is_table_61 AND is_central_pcs;
	wire_w_lg_is_tier_1246w(0) <= is_tier_1 AND wire_w_lg_header_proc225w(0);
	wire_w_lg_is_tier_1221w(0) <= is_tier_1 AND wire_w_lg_w219w220w(0);
	wire_w_lg_is_tier_1206w(0) <= is_tier_1 AND mif_reconfig_done;
	wire_w_lg_read49w(0) <= read AND en_read_trigger;
	loop13 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_read_address192w(i) <= read_address(i) AND read_state;
	END GENERATE loop13;
	wire_w_lg_read_state214w(0) <= read_state AND wire_w_lg_dprio_pulse213w(0);
	wire_w_lg_read_state727w(0) <= read_state AND read_word_7c_7f_data_valid;
	loop14 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state681w(i) <= read_state AND w_rx_eqctrl_out567w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_read_state701w(i) <= read_state AND w_rx_eqdcgain_out683w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_read_state724w(i) <= read_state AND w_tx_vodctrl_out703w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_read_state737w(i) <= read_state AND wire_dprio_w_dataout_range410w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state731w(i) <= read_state AND wire_dprio_w_dataout_range730w(i);
	END GENERATE loop18;
	wire_w_lg_read_state760w(0) <= read_state AND wire_dprio_w_dataout_range759w(0);
	wire_w_lg_read_state750w(0) <= read_state AND wire_dprio_w_dataout_range749w(0);
	loop19 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state743w(i) <= read_state AND wire_dprio_w_dataout_range742w(i);
	END GENERATE loop19;
	wire_w_lg_read_word_64_67_data_valid698w(0) <= read_word_64_67_data_valid AND read_state;
	wire_w_lg_read_word_68_6B_data_valid678w(0) <= read_word_68_6B_data_valid AND read_state;
	wire_w_lg_read_word_7c_7f_data_valid739w(0) <= read_word_7c_7f_data_valid AND read_state;
	wire_w_lg_read_word_7c_7f_inv_data_valid316w(0) <= read_word_7c_7f_inv_data_valid AND wire_w_lg_rx_reconfig315w(0);
	wire_w_lg_read_word_preemp_1t_data_valid734w(0) <= read_word_preemp_1t_data_valid AND read_state;
	wire_w_lg_read_word_vodctrl_data_valid721w(0) <= read_word_vodctrl_data_valid AND read_state;
	loop20 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_0_617w673w(i) <= w_eq_0_617w(i) AND w_gt_0_only601w;
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_10_658w670w(i) <= w_eq_10_658w(i) AND w_gt_10_only615w;
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_3_639w672w(i) <= w_eq_3_639w(i) AND w_gt_3_only608w;
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_6_649w671w(i) <= w_eq_6_649w(i) AND w_gt_6_only612w;
	END GENERATE loop23;
	wire_w_lg_w_gt_0_577w605w(0) <= w_gt_0_577w AND wire_w_lg_w_gt_3_583w604w(0);
	wire_w_lg_w_gt_0_577w609w(0) <= w_gt_0_577w AND w_gt_3_583w;
	wire_w_lg_wr_pulse345w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q337w(0);
	wire_w_lg_wr_pulse342w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q341w(0);
	loop24 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_address193w(i) <= write_address(i) AND write_state;
	END GENERATE loop24;
	wire_w_lg_write_all25w(0) <= write_all AND wire_w_lg_w_lg_is_bonded_reconfig17w24w(0);
	wire_w_lg_write_state228w(0) <= write_state AND wire_w_lg_w_lg_w_lg_header_proc225w226w227w(0);
	wire_w_lg_write_state252w(0) <= write_state AND wire_w_lg_dprio_pulse213w(0);
	wire_w_lg_write_state748w(0) <= write_state AND wire_w_lg_w_tx_preemp_0t_range2w509w(0);
	wire_w_lg_write_state758w(0) <= write_state AND wire_w_lg_w_tx_preemp_2t_range4w513w(0);
	loop25 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state680w(i) <= write_state AND rx_eqctrl(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_state700w(i) <= write_state AND rx_eqdcgain(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_write_state736w(i) <= write_state AND tx_preemp_1t(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_state723w(i) <= write_state AND tx_vodctrl(i);
	END GENERATE loop28;
	wire_w_lg_write_state697w(0) <= write_state AND write_word_64_67_data_valid;
	wire_w_lg_write_state677w(0) <= write_state AND write_word_68_6B_data_valid;
	wire_w_lg_write_state726w(0) <= write_state AND write_word_7c_7f_data_valid;
	wire_w_lg_write_state733w(0) <= write_state AND write_word_preemp1t_data_valid;
	wire_w_lg_write_state720w(0) <= write_state AND write_word_vodctrl_data_valid;
	loop29 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state729w(i) <= write_state AND wire_w_tx_preemp_0t_wire_range507w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state741w(i) <= write_state AND wire_w_tx_preemp_2t_wire_range511w(i);
	END GENERATE loop30;
	wire_w_lg_write_word_7c_7f_inv_data_valid551w(0) <= write_word_7c_7f_inv_data_valid AND wire_w_lg_rx_reconfig315w(0);
	wire_w_lg_write_word_done519w(0) <= write_word_done AND write_addr_inc;
	wire_w_lg_w_rx_eqctrl_range451w467w(0) <= wire_w_rx_eqctrl_range451w(0) AND wire_w_lg_w_rx_eqctrl_range458w466w(0);
	wire_w_lg_w_rx_eqctrl_range451w477w(0) <= wire_w_rx_eqctrl_range451w(0) AND wire_w_lg_w_rx_eqctrl_range458w476w(0);
	wire_w_lg_w_rx_eqctrl_range453w461w(0) <= wire_w_rx_eqctrl_range453w(0) AND wire_w_lg_w_rx_eqctrl_range451w452w(0);
	wire_w_lg_w_rx_eqctrl_range453w484w(0) <= wire_w_rx_eqctrl_range453w(0) AND wire_w_rx_eqctrl_range451w(0);
	wire_w_lg_w_rx_eqctrl_range455w456w(0) <= wire_w_rx_eqctrl_range455w(0) AND wire_w_lg_w_rx_eqctrl_range453w454w(0);
	wire_w_lg_w_rx_eqctrl_range455w482w(0) <= wire_w_rx_eqctrl_range455w(0) AND wire_w_rx_eqctrl_range451w(0);
	wire_w_lg_w_rx_eqctrl_range455w459w(0) <= wire_w_rx_eqctrl_range455w(0) AND wire_w_rx_eqctrl_range453w(0);
	wire_w_lg_w_rx_eqdcgain_range433w434w(0) <= wire_w_rx_eqdcgain_range433w(0) AND wire_w_rx_eqdcgain_range432w(0);
	wire_w_lg_w_tx_vodctrl_range374w382w(0) <= wire_w_tx_vodctrl_range374w(0) AND wire_w_lg_w_lg_w_tx_vodctrl_range372w373w381w(0);
	wire_w_lg_w_tx_vodctrl_range374w375w(0) <= wire_w_tx_vodctrl_range374w(0) AND wire_w_lg_w_tx_vodctrl_range372w373w(0);
	wire_w_lg_w_tx_vodctrl_range372w384w(0) <= wire_w_tx_vodctrl_range372w(0) AND wire_w_lg_w_tx_vodctrl_range371w383w(0);
	wire_w_lg_w_tx_vodctrl_range372w376w(0) <= wire_w_tx_vodctrl_range372w(0) AND wire_w_tx_vodctrl_range371w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w628w(0) <= wire_w_w_rx_eqv572w_range627w(0) AND wire_w_lg_w_lg_w_w_rx_eqv572w_range624w625w626w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w646w(0) <= wire_w_w_rx_eqv572w_range627w(0) AND wire_w_lg_w_w_rx_eqv572w_range624w631w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w635w(0) <= wire_w_w_rx_eqv572w_range627w(0) AND wire_w_w_rx_eqv572w_range624w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range455w486w487w(0) <= NOT wire_w_lg_w_rx_eqctrl_range455w486w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range372w373w381w(0) <= NOT wire_w_lg_w_tx_vodctrl_range372w373w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range624w625w626w(0) <= NOT wire_w_lg_w_w_rx_eqv572w_range624w625w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range627w654w655w(0) <= NOT wire_w_lg_w_w_rx_eqv572w_range627w654w(0);
	wire_w_lg_bonded_skip237w(0) <= NOT bonded_skip;
	wire_w_lg_cal_busy89w(0) <= NOT cal_busy;
	wire_w_lg_dprio_pulse213w(0) <= NOT dprio_pulse;
	wire_w_lg_header_proc225w(0) <= NOT header_proc;
	wire_w_lg_is_analog_control344w(0) <= NOT is_analog_control;
	wire_w_lg_is_bonded_global_clk_div9w(0) <= NOT is_bonded_global_clk_div;
	wire_w_lg_is_bonded_reconfig17w(0) <= NOT is_bonded_reconfig;
	wire_w_lg_is_central_pcs118w(0) <= NOT is_central_pcs;
	wire_w_lg_is_cruclk_addr0239w(0) <= NOT is_cruclk_addr0;
	wire_w_lg_is_diff_mif196w(0) <= NOT is_diff_mif;
	wire_w_lg_is_global_clk_div_mode235w(0) <= NOT is_global_clk_div_mode;
	wire_w_lg_is_illegal_reg_d211w(0) <= NOT is_illegal_reg_d;
	wire_w_lg_is_pll_address106w(0) <= NOT is_pll_address;
	wire_w_lg_is_protected_bit236w(0) <= NOT is_protected_bit;
	wire_w_lg_is_rcxpat_chnl_en_ch240w(0) <= NOT is_rcxpat_chnl_en_ch;
	wire_w_lg_is_table_3313w(0) <= NOT is_table_33;
	wire_w_lg_is_tier_1222w(0) <= NOT is_tier_1;
	wire_w_lg_rd_pulse143w(0) <= NOT rd_pulse;
	wire_w_lg_read_done212w(0) <= NOT read_done;
	wire_w_lg_read_state203w(0) <= NOT read_state;
	wire_w_lg_reset_reconf_addr224w(0) <= NOT reset_reconf_addr;
	wire_w_lg_rx_reconfig315w(0) <= NOT rx_reconfig;
	wire_w_lg_s0_to_056w(0) <= NOT s0_to_0;
	wire_w_lg_s0_to_157w(0) <= NOT s0_to_1;
	wire_w_lg_s1_to_068w(0) <= NOT s1_to_0;
	wire_w_lg_s1_to_169w(0) <= NOT s1_to_1;
	wire_w_lg_s2_to_058w(0) <= NOT s2_to_0;
	wire_w_lg_tx_reconfig294w(0) <= NOT tx_reconfig;
	wire_w_lg_w_gt_10_595w602w(0) <= NOT w_gt_10_595w;
	wire_w_lg_w_gt_3_583w604w(0) <= NOT w_gt_3_583w;
	wire_w_lg_w_gt_6_589w603w(0) <= NOT w_gt_6_589w;
	wire_w_lg_wr_pulse144w(0) <= NOT wr_pulse;
	wire_w_lg_write_all_int47w(0) <= NOT write_all_int;
	wire_w_lg_write_done229w(0) <= NOT write_done;
	wire_w_lg_write_skip238w(0) <= NOT write_skip;
	wire_w_lg_write_state48w(0) <= NOT write_state;
	wire_w_lg_w_reconfig_mode_sel_range76w77w(0) <= NOT wire_w_reconfig_mode_sel_range76w(0);
	wire_w_lg_w_reconfig_mode_sel_range81w82w(0) <= NOT wire_w_reconfig_mode_sel_range81w(0);
	wire_w_lg_w_rx_eqctrl_range458w466w(0) <= NOT wire_w_rx_eqctrl_range458w(0);
	wire_w_lg_w_rx_eqctrl_range451w452w(0) <= NOT wire_w_rx_eqctrl_range451w(0);
	wire_w_lg_w_rx_eqctrl_range453w454w(0) <= NOT wire_w_rx_eqctrl_range453w(0);
	wire_w_lg_w_rx_eqctrl_range455w463w(0) <= NOT wire_w_rx_eqctrl_range455w(0);
	wire_w_lg_w_tx_preemp_0t_range2w509w(0) <= NOT wire_w_tx_preemp_0t_range2w(0);
	wire_w_lg_w_tx_preemp_2t_range4w513w(0) <= NOT wire_w_tx_preemp_2t_range4w(0);
	wire_w_lg_w_tx_vodctrl_range371w383w(0) <= NOT wire_w_tx_vodctrl_range371w(0);
	wire_w_lg_w_w_rx_eqv572w_range623w630w(0) <= NOT wire_w_w_rx_eqv572w_range623w(0);
	wire_w_lg_w_w_rx_eqv572w_range624w631w(0) <= NOT wire_w_w_rx_eqv572w_range624w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w632w(0) <= NOT wire_w_w_rx_eqv572w_range627w(0);
	wire_w_lg_w489w490w(0) <= wire_w489w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range453w484w485w(0);
	wire_w637w(0) <= wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w(0) OR wire_w634w(0);
	wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w(0) <= wire_w_lg_w_lg_is_bonded_global_clk_div9w10w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_w_lg_is_table_3313w14w15w(0) <= wire_w_lg_w_lg_is_table_3313w14w(0) OR wire_w_lg_is_table_3312w(0);
	wire_w665w(0) <= wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w656w(0) OR wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w(0);
	wire_w668w(0) <= wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w667w(0) OR wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w(0);
	wire_w_lg_w_lg_w125w126w127w(0) <= wire_w_lg_w125w126w(0) OR wire_w_lg_is_table_61117w(0);
	wire_w125w(0) <= wire_w_lg_w_lg_w_channel_address_range122w123w124w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range119w120w121w(0);
	wire_w110w(0) <= wire_w_lg_w_lg_w_channel_address_range107w108w109w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range103w104w105w(0);
	loop31 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_cal_busy91w92w(i) <= wire_w_lg_cal_busy91w(i) OR wire_w_lg_w_lg_cal_busy89w90w(i);
	END GENERATE loop31;
	wire_w_lg_w_lg_cal_busy130w131w(0) <= wire_w_lg_cal_busy130w(0) OR wire_w_lg_w_lg_cal_busy89w128w(0);
	wire_w_lg_w_lg_cal_busy114w115w(0) <= wire_w_lg_cal_busy114w(0) OR wire_w_lg_w_lg_cal_busy89w112w(0);
	wire_w_lg_w_lg_cal_busy99w100w(0) <= wire_w_lg_cal_busy99w(0) OR wire_w_lg_w_lg_cal_busy89w97w(0);
	loop32 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_vodctrl362w363w(i) <= wire_w_lg_dprio_datain_vodctrl362w(i) OR wire_w_lg_dprio_datain_preemp1t360w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_read_state727w728w(0) <= wire_w_lg_read_state727w(0) OR wire_w_lg_write_state726w(0);
	loop33 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state681w682w(i) <= wire_w_lg_read_state681w(i) OR wire_w_lg_write_state680w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_read_state701w702w(i) <= wire_w_lg_read_state701w(i) OR wire_w_lg_write_state700w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_read_state724w725w(i) <= wire_w_lg_read_state724w(i) OR wire_w_lg_write_state723w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_read_state737w738w(i) <= wire_w_lg_read_state737w(i) OR wire_w_lg_write_state736w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state731w732w(i) <= wire_w_lg_read_state731w(i) OR wire_w_lg_write_state729w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state743w744w(i) <= wire_w_lg_read_state743w(i) OR wire_w_lg_write_state741w(i);
	END GENERATE loop38;
	wire_w_lg_w_lg_read_word_64_67_data_valid698w699w(0) <= wire_w_lg_read_word_64_67_data_valid698w(0) OR wire_w_lg_write_state697w(0);
	wire_w_lg_w_lg_read_word_68_6B_data_valid678w679w(0) <= wire_w_lg_read_word_68_6B_data_valid678w(0) OR wire_w_lg_write_state677w(0);
	wire_w_lg_w_lg_read_word_7c_7f_data_valid739w740w(0) <= wire_w_lg_read_word_7c_7f_data_valid739w(0) OR wire_w_lg_write_state726w(0);
	wire_w_lg_w_lg_read_word_preemp_1t_data_valid734w735w(0) <= wire_w_lg_read_word_preemp_1t_data_valid734w(0) OR wire_w_lg_write_state733w(0);
	wire_w_lg_w_lg_read_word_vodctrl_data_valid721w722w(0) <= wire_w_lg_read_word_vodctrl_data_valid721w(0) OR wire_w_lg_write_state720w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range451w467w468w(0) <= wire_w_lg_w_rx_eqctrl_range451w467w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w463w464w465w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range451w477w478w(0) <= wire_w_lg_w_rx_eqctrl_range451w477w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w459w473w474w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range372w384w385w(0) <= wire_w_lg_w_tx_vodctrl_range372w384w(0) OR wire_w_lg_w_tx_vodctrl_range374w382w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range372w376w377w(0) <= wire_w_lg_w_tx_vodctrl_range372w376w(0) OR wire_w_lg_w_tx_vodctrl_range374w375w(0);
	wire_w_lg_w_lg_is_bonded_reconfig17w24w(0) <= wire_w_lg_is_bonded_reconfig17w(0) OR wire_w_lg_is_bonded_reconfig23w(0);
	wire_w_lg_w_lg_is_tier_1222w249w(0) <= wire_w_lg_is_tier_1222w(0) OR wire_w_lg_w_lg_is_tier_1246w248w(0);
	wire_w_lg_w_lg_is_tier_1222w223w(0) <= wire_w_lg_is_tier_1222w(0) OR wire_w_lg_is_tier_1221w(0);
	wire_w_lg_w_lg_w489w490w491w(0) <= wire_w_lg_w489w490w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range455w482w483w(0);
	wire_w_lg_w110w111w(0) <= wire_w110w(0) OR is_central_pcs;
	loop39 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl362w363w364w(i) <= wire_w_lg_w_lg_dprio_datain_vodctrl362w363w(i) OR wire_w_lg_dprio_datain_64_67357w(i);
	END GENERATE loop39;
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range451w467w468w469w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range451w467w468w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range453w461w462w(0);
	wire_w_lg_w_lg_w_lg_w489w490w491w492w(0) <= wire_w_lg_w_lg_w489w490w491w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range455w459w481w(0);
	loop40 : FOR i IN 0 TO 15 GENERATE 
		wire_w365w(i) <= wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl362w363w364w(i) OR wire_w_lg_w_lg_dprio_datain_68_6B355w356w(i);
	END GENERATE loop40;
	wire_w470w(0) <= wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range451w467w468w469w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range455w459w460w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w489w490w491w492w493w(0) <= wire_w_lg_w_lg_w_lg_w489w490w491w492w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range455w456w457w480w(0);
	loop41 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w365w366w(i) <= wire_w365w(i) OR wire_w_lg_dprio_datain_7c_7f354w(i);
	END GENERATE loop41;
	wire_w_lg_w470w471w(0) <= wire_w470w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range455w456w457w(0);
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w365w366w367w(i) <= wire_w_lg_w365w366w(i) OR wire_w_lg_dprio_datain_7c_7f_inv353w(i);
	END GENERATE loop42;
	wire_w_lg_w219w220w(0) <= wire_w219w(0) OR is_global_clk_div_mode;
	wire_w219w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w218w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w218w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w(0) OR bonded_skip;
	wire_w_lg_w_lg_is_adce39w40w(0) <= wire_w_lg_is_adce39w(0) OR is_do_dfe;
	wire_w_lg_w_lg_is_pll_address95w96w(0) <= wire_w_lg_is_pll_address95w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch216w217w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch216w(0) OR write_skip;
	wire_w_lg_w_lg_is_tier_1350w351w(0) <= wire_w_lg_is_tier_1350w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_s0_to_262w63w(0) <= wire_w_lg_s0_to_262w(0) OR wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w(0);
	wire_w_lg_w_lg_s0_to_273w74w(0) <= wire_w_lg_s0_to_273w(0) OR wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w(0);
	wire_w_lg_w_lg_write_word_preemp1t_data_valid358w359w(0) <= wire_w_lg_write_word_preemp1t_data_valid358w(0) OR write_word_preemp1tb_data_valid;
	wire_w_lg_w_lg_w_rx_eqdcgain_range429w437w439w(0) <= wire_w_lg_w_rx_eqdcgain_range429w437w(0) OR wire_w_rx_eqdcgain_range432w(0);
	wire_w_lg_w_lg_w_w_rx_eqv572w_range627w662w663w(0) <= wire_w_lg_w_w_rx_eqv572w_range627w662w(0) OR wire_w_w_rx_eqv572w_range623w(0);
	loop43 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_68_6B355w(i) <= dprio_datain_68_6B(i) OR local_ch_dec;
	END GENERATE loop43;
	wire_w_lg_is_adce39w(0) <= is_adce OR is_do_eyemon;
	wire_w_lg_is_pll_address95w(0) <= is_pll_address OR is_central_pcs;
	wire_w_lg_is_rcxpat_chnl_en_ch216w(0) <= is_rcxpat_chnl_en_ch OR is_cruclk_addr0;
	wire_w_lg_is_tier_1350w(0) <= is_tier_1 OR is_tier_2;
	wire_w_lg_reset_system207w(0) <= reset_system OR wire_w_lg_is_tier_1206w(0);
	wire_w_lg_s0_to_262w(0) <= s0_to_2 OR s0_to_1;
	wire_w_lg_s0_to_273w(0) <= s0_to_2 OR s1_to_1;
	wire_w_lg_write_word_preemp1t_data_valid358w(0) <= write_word_preemp1t_data_valid OR write_word_preemp1ta_data_valid;
	wire_w_lg_write_word_vodctrl_data_valid361w(0) <= write_word_vodctrl_data_valid OR write_word_vodctrla_data_valid;
	wire_w_lg_w_channel_address_range122w123w(0) <= wire_w_channel_address_range122w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_channel_address_range107w108w(0) <= wire_w_channel_address_range107w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_logical_pll_sel_num_range119w120w(0) <= wire_w_logical_pll_sel_num_range119w(0) OR wire_w_lg_is_table_59102w(0);
	wire_w_lg_w_logical_pll_sel_num_range103w104w(0) <= wire_w_logical_pll_sel_num_range103w(0) OR wire_w_lg_is_table_59102w(0);
	wire_w_lg_w_reconfig_mode_sel_range81w87w(0) <= wire_w_reconfig_mode_sel_range81w(0) OR wire_w86w(0);
	wire_w_lg_w_rx_eqdcgain_range429w435w(0) <= wire_w_rx_eqdcgain_range429w(0) OR wire_w_lg_w_rx_eqdcgain_range433w434w(0);
	wire_w_lg_w_rx_eqdcgain_range429w437w(0) <= wire_w_rx_eqdcgain_range429w(0) OR wire_w_rx_eqdcgain_range433w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w662w(0) <= wire_w_w_rx_eqv572w_range627w(0) OR wire_w_w_rx_eqv572w_range624w(0);
	wire_w_lg_w_rx_eqctrl_range458w476w(0) <= wire_w_rx_eqctrl_range458w(0) XOR wire_w_lg_w_rx_eqctrl_range453w475w(0);
	wire_w_lg_w_rx_eqctrl_range453w475w(0) <= wire_w_rx_eqctrl_range453w(0) XOR wire_w_rx_eqctrl_range455w(0);
	wire_w_lg_w_rx_eqctrl_range455w486w(0) <= wire_w_rx_eqctrl_range455w(0) XOR wire_w_rx_eqctrl_range453w(0);
	wire_w_lg_w_tx_vodctrl_range372w373w(0) <= wire_w_tx_vodctrl_range372w(0) XOR wire_w_tx_vodctrl_range371w(0);
	wire_w_lg_w_w_rx_eqv572w_range624w625w(0) <= wire_w_w_rx_eqv572w_range624w(0) XOR wire_w_w_rx_eqv572w_range623w(0);
	wire_w_lg_w_w_rx_eqv572w_range627w654w(0) <= wire_w_w_rx_eqv572w_range627w(0) XOR wire_w_w_rx_eqv572w_range623w(0);
	a2gr_dprio_addr <= (wire_w_lg_write_address193w OR wire_w_lg_read_address192w);
	a2gr_dprio_data <= wire_w_lg_w_lg_dprio_datain348w349w;
	a2gr_dprio_rden <= (rd_pulse AND (wire_w_lg_is_diff_mif196w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren <= ((wire_w_lg_wr_pulse345w(0) AND wire_w_lg_is_analog_control344w(0)) AND (wire_w_lg_is_diff_mif196w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren_data <= (wire_w_lg_wr_pulse342w(0) AND (wire_w_lg_is_diff_mif196w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	adce_busy_state <= '0';
	adce_state <= (state_mc_reg(0) AND state_mc_reg(1));
	aeq_ch_done <= (OTHERS => '0');
	bonded_skip <= '0';
	busy <= (((wire_w_lg_w_lg_is_bonded_reconfig17w18w(0) OR wire_w_lg_is_bonded_reconfig16w(0)) OR internal_write_pulse) OR cal_busy);
	busy_state <= ((((read_state OR write_state) OR adce_state) OR eyemon_busy) OR dfe_busy);
	cal_busy <= wire_calibration_busy;
	cal_channel_address <= wire_calibration_dprio_addr(14 DOWNTO 12);
	cal_channel_address_out <= address_pres_reg(2 DOWNTO 0);
	cal_dprio_address <= ( wire_calibration_dprio_addr(15) & cal_channel_address_out & wire_calibration_dprio_addr(11 DOWNTO 0));
	cal_dprioout_wire <= ( reconfig_fromgxb(17) & reconfig_fromgxb(0));
	cal_quad_address <= wire_calibration_quad_addr;
	cal_testbuses <= ( reconfig_fromgxb(33 DOWNTO 18) & reconfig_fromgxb(16 DOWNTO 1));
	channel_address <= wire_addr_cntr_q(1 DOWNTO 0);
	channel_address_out <= wire_address_pres_reg_w_lg_w_q_range140w141w;
	data_valid <= (data_valid_reg AND idle_state);
	dfe_busy <= '0';
	diff_mif_wr_rd_busy <= '0';
	dprio_datain <= (wire_w_lg_w_lg_w_lg_w365w366w367w368w OR wire_w_lg_w_lg_w_lg_is_tier_1350w351w352w);
	dprio_datain_64_67 <= ( wire_dprio_dataout(15 DOWNTO 11) & ( rx_eqdcgain(2) & wire_w_lg_w_rx_eqdcgain_range429w435w & wire_w_lg_w_rx_eqdcgain_range429w437w & wire_w_lg_w_lg_w_rx_eqdcgain_range429w437w439w) & wire_dprio_dataout(6 DOWNTO 0));
	dprio_datain_68_6B <= ( wire_dprio_dataout(15) & ( wire_cmpr6_agb & wire_cmpr6_agb & wire_cmpr6_agb & wire_cmpr7_agb & wire_cmpr7_agb & wire_cmpr7_agb & wire_cmpr8_agb & wire_cmpr8_agb & wire_cmpr8_agb & wire_cmpr9_agb & wire_cmpr9_agb & wire_cmpr9_agb & wire_w_lg_w470w471w & wire_w_lg_w_lg_w_rx_eqctrl_range451w477w478w & wire_w_lg_w_lg_w_lg_w_lg_w489w490w491w492w493w));
	dprio_datain_7c_7f <= ( wire_dprio_dataout(15 DOWNTO 8) & tx_preemp_2t_wire(3 DOWNTO 0) & tx_preemp_0t_wire(3 DOWNTO 0));
	dprio_datain_7c_7f_inv <= ( wire_dprio_dataout(15 DOWNTO 5) & wire_w_lg_w_tx_preemp_0t_range2w509w & wire_w_lg_w_tx_preemp_2t_range4w513w & wire_dprio_dataout(2 DOWNTO 0));
	dprio_datain_preemp1t <= ( tx_preemp_1t & wire_dprio_dataout(10 DOWNTO 0));
	dprio_datain_vodctrl <= ( ( wire_w_lg_w_lg_w_tx_vodctrl_range372w376w377w & wire_w_lg_w_tx_vodctrl_range372w373w & wire_w_lg_w_lg_w_tx_vodctrl_range372w384w385w) & wire_dprio_dataout(12 DOWNTO 0));
	dprio_pulse <= ((dprio_pulse_reg XOR wire_dprio_busy) AND wire_dprio_w_lg_busy199w(0));
	en_read_trigger <= legal_rd_mode_type;
	en_write_trigger <= legal_wr_mode_type;
	eyemon_busy <= '0';
	header_proc <= '0';
	idle_state <= (wire_state_mc_reg_w_lg_q31w(0) AND wire_state_mc_reg_w_lg_q29w(0));
	internal_write_pulse <= '0';
	is_adce <= ((((is_adce_single_control OR is_adce_all_control) OR is_adce_continuous_single_control) OR is_adce_one_time_single_control) OR is_adce_standby_single_control);
	is_adce_all_control <= '0';
	is_adce_continuous_single_control <= '0';
	is_adce_one_time_single_control <= '0';
	is_adce_single_control <= '0';
	is_adce_standby_single_control <= '0';
	is_analog_control <= wire_reconf_mode_dec_eq(0);
	is_bonded_global_clk_div <= '0';
	is_bonded_reconfig <= '0';
	is_central_pcs <= '0';
	is_cruclk_addr0 <= '0';
	is_diff_mif <= '0';
	is_do_dfe <= '0';
	is_do_eyemon <= '0';
	is_illegal_reg_d <= '0';
	is_illegal_reg_out <= '0';
	is_pll_address <= '0';
	is_protected_bit <= '0';
	is_rcxpat_chnl_en_ch <= '0';
	is_table_33 <= '0';
	is_table_59 <= '0';
	is_table_61 <= '0';
	is_tier_1 <= '0';
	is_tier_2 <= '0';
	is_tx_local_div_ctrl <= '0';
	legal_rd_mode_type <= (wire_w_lg_w_reconfig_mode_sel_range81w82w(0) AND ((NOT reconfig_mode_sel(1)) AND wire_w_lg_w_reconfig_mode_sel_range76w77w(0)));
	legal_wr_mode_type <= (wire_w_lg_w_reconfig_mode_sel_range81w87w(0) OR (wire_w_lg_w_reconfig_mode_sel_range81w82w(0) AND (NOT reconfig_mode_sel(1))));
	local_ch_dec <= wire_aeq_ch_done_mux_result(0);
	logical_pll_sel_num <= (OTHERS => '0');
	mif_reconfig_done <= '0';
	quad_address <= ( "00000000" & wire_addr_cntr_q(2));
	quad_address_out <= address_pres_reg(11 DOWNTO 3);
	rd_pulse <= (((((wire_w_lg_dprio_pulse213w(0) AND wire_w_lg_write_done229w(0)) AND wire_wr_rd_pulse_reg_w_lg_q202w(0)) AND wire_w_lg_write_state228w(0)) OR (wire_w_lg_read_state214w(0) AND wire_w_lg_read_done212w(0))) AND wire_w_lg_is_illegal_reg_d211w(0));
	read_addr_inc <= (read_state AND dprio_pulse);
	read_address <= ( "0" & address_pres_reg(2) & channel_address_out & "1" & wire_read_addr_cntr_q(2) & "000000" & wire_read_addr_cntr_w_lg_w_q_range305w308w & "0" & wire_read_addr_cntr_w_lg_w_q_range311w312w & wire_read_addr_cntr_q(0));
	read_done <= (((read_word_done AND read_addr_inc) OR (is_illegal_reg_out AND read_state)) OR reset_system);
	read_state <= (state_mc_reg(0) AND wire_state_mc_reg_w_lg_q29w(0));
	read_word_64_67_data_valid <= ((wire_w_lg_dprio_pulse329w(0) AND (NOT wire_read_addr_cntr_q(1))) AND (NOT wire_read_addr_cntr_q(0)));
	read_word_68_6B_data_valid <= ((wire_w_lg_dprio_pulse329w(0) AND (NOT wire_read_addr_cntr_q(1))) AND wire_read_addr_cntr_q(0));
	read_word_7c_7f_data_valid <= ((wire_w_lg_dprio_pulse322w(0) AND wire_read_addr_cntr_q(1)) AND (NOT wire_read_addr_cntr_q(0)));
	read_word_7c_7f_inv_data_valid <= ((wire_w_lg_dprio_pulse322w(0) AND wire_read_addr_cntr_q(1)) AND wire_read_addr_cntr_q(0));
	read_word_done <= ((read_word_68_6B_data_valid AND rx_reconfig) OR wire_w_lg_read_word_7c_7f_inv_data_valid316w(0));
	read_word_preemp_1t_data_valid <= ((wire_w_lg_dprio_pulse322w(0) AND (NOT wire_read_addr_cntr_q(1))) AND wire_read_addr_cntr_q(0));
	read_word_vodctrl_data_valid <= ((wire_w_lg_dprio_pulse322w(0) AND (NOT wire_read_addr_cntr_q(1))) AND (NOT wire_read_addr_cntr_q(0)));
	reconfig_datain <= (OTHERS => '0');
	reconfig_reset_all <= '0';
	reconfig_togxb <= ( wire_calibration_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	reset_addr_done <= '0';
	reset_reconf_addr <= '0';
	reset_system <= '0';
	rx_eqctrl_out <= rx_eqctrl_reg;
	rx_eqdcgain_out <= rx_equalizer_dcgain_reg;
	rx_reconfig <= '1';
	s0_to_0 <= ((idle_state AND write_all_int) OR read_done);
	s0_to_1 <= ((wire_w_lg_idle_state50w(0) AND wire_w_lg_write_state48w(0)) AND wire_w_lg_write_all_int47w(0));
	s0_to_2 <= (wire_w_lg_idle_state41w(0) AND (wire_w_lg_write_all25w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)));
	s1_to_0 <= ((wire_w_lg_idle_state50w(0) AND wire_w_lg_write_state48w(0)) OR write_done);
	s1_to_1 <= (idle_state AND write_all_int);
	s2_to_0 <= (adce_state AND (NOT ((adce_busy_state OR eyemon_busy) OR dfe_busy)));
	start <= '0';
	state_mc_reg_in <= ( wire_w_lg_w_lg_s0_to_273w74w & wire_w_lg_w_lg_s0_to_262w63w);
	transceiver_init <= '0';
	tx_preemp_0t_out <= ( wire_tx_preemp_0t_inv_reg_w_lg_w_q_range752w753w & wire_add_sub10_result);
	tx_preemp_0t_out_wire <= tx_preemphasisctrl_pretap_reg;
	tx_preemp_0t_wire <= wire_add_sub1_result;
	tx_preemp_1t_out <= tx_preemphasisctrl_1stposttap_reg;
	tx_preemp_2t_out <= ( wire_tx_preemp_2t_inv_reg_w_lg_w_q_range762w763w & wire_add_sub11_result);
	tx_preemp_2t_out_wire <= tx_preemphasisctrl_2ndposttap_reg;
	tx_preemp_2t_wire <= wire_add_sub2_result;
	tx_reconfig <= '1';
	tx_vodctrl_out <= tx_vodctrl_reg;
	w334w <= ( quad_address & channel_address);
	w_eq_0_617w <= ( "0" & "0" & wire_w_lg_w_w_rx_eqv572w_range627w628w & wire_w637w);
	w_eq_10_658w <= ( "1" & wire_w_lg_w_lg_w_w_rx_eqv572w_range627w662w663w & wire_w665w & wire_w668w);
	w_eq_3_639w <= ( "0" & "1" & wire_w_lg_w_lg_w_w_rx_eqv572w_range627w635w636w & wire_w_lg_w_lg_w_w_rx_eqv572w_range627w646w647w);
	w_eq_6_649w <= ( w_rx_eqv572w(2) & wire_w_lg_w_w_rx_eqv572w_range627w632w & wire_w637w & wire_w_lg_w_lg_w_w_rx_eqv572w_range624w631w656w);
	w_gt_0_577w <= ((w_rx_eqd568w(2) AND w_rx_eqd568w(1)) AND w_rx_eqd568w(0));
	w_gt_0_only601w <= ((wire_w_lg_w_gt_0_577w605w(0) AND wire_w_lg_w_gt_6_589w603w(0)) AND wire_w_lg_w_gt_10_595w602w(0));
	w_gt_10_595w <= ((w_rx_eqa571w(2) AND w_rx_eqa571w(1)) AND w_rx_eqa571w(0));
	w_gt_10_only615w <= (wire_w_lg_w_lg_w_gt_0_577w609w613w(0) AND ((w_rx_eqa571w(2) AND w_rx_eqa571w(1)) AND w_rx_eqa571w(0)));
	w_gt_3_583w <= ((w_rx_eqc569w(2) AND w_rx_eqc569w(1)) AND w_rx_eqc569w(0));
	w_gt_3_only608w <= ((wire_w_lg_w_gt_0_577w609w(0) AND wire_w_lg_w_gt_6_589w603w(0)) AND wire_w_lg_w_gt_10_595w602w(0));
	w_gt_6_589w <= ((w_rx_eqb570w(2) AND w_rx_eqb570w(1)) AND w_rx_eqb570w(0));
	w_gt_6_only612w <= (wire_w_lg_w_lg_w_gt_0_577w609w613w(0) AND wire_w_lg_w_gt_10_595w602w(0));
	w_rx_eqa571w <= wire_dprio_dataout(14 DOWNTO 12);
	w_rx_eqb570w <= wire_dprio_dataout(11 DOWNTO 9);
	w_rx_eqc569w <= wire_dprio_dataout(8 DOWNTO 6);
	w_rx_eqctrl_out567w <= (((wire_w_lg_w_eq_0_617w673w OR wire_w_lg_w_eq_3_639w672w) OR wire_w_lg_w_eq_6_649w671w) OR wire_w_lg_w_eq_10_658w670w);
	w_rx_eqd568w <= wire_dprio_dataout(5 DOWNTO 3);
	w_rx_eqdcgain_out683w <= ( wire_dprio_dataout(10) & wire_dprio_w_lg_w_dataout_range688w689w & wire_dprio_w_lg_w_lg_w_lg_w_dataout_range692w693w694w695w);
	w_rx_eqv572w <= wire_dprio_dataout(2 DOWNTO 0);
	w_tx_vodctrl_out703w <= ( wire_dprio_w_lg_w_lg_w_dataout_range704w708w709w & wire_dprio_w_lg_w_lg_w_dataout_range704w713w714w & wire_dprio_w_lg_w_lg_w_lg_w_dataout_range704w705w717w718w);
	wr_pulse <= (((wire_w_lg_write_state252w(0) AND wire_w_lg_write_done229w(0)) AND (wire_wr_rd_pulse_reg_w_lg_q250w(0) OR (wire_w_lg_is_tier_1246w(0) AND (((((wire_w_lg_is_rcxpat_chnl_en_ch240w(0) AND wire_w_lg_is_cruclk_addr0239w(0)) AND wire_w_lg_write_skip238w(0)) AND wire_w_lg_bonded_skip237w(0)) AND wire_w_lg_is_protected_bit236w(0)) AND wire_w_lg_is_global_clk_div_mode235w(0))))) AND wire_w_lg_is_illegal_reg_d211w(0));
	write_addr_inc <= ((write_state AND dprio_pulse) AND write_happened);
	write_address <= ( "0" & address_pres_reg(2) & channel_address_out & "1" & wire_write_addr_cntr_q(2) & "000000" & wire_write_addr_cntr_w_lg_w_q_range541w544w & "0" & wire_write_addr_cntr_w_lg_w_q_range547w548w & wire_write_addr_cntr_q(0));
	write_all_int <= ((wire_w_lg_write_all25w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)) AND en_write_trigger);
	write_done <= ((wire_w_lg_w_lg_write_word_done519w520w(0) OR (is_illegal_reg_out AND write_state)) OR reset_system);
	write_happened <= wr_addr_inc_reg;
	write_skip <= '0';
	write_state <= (wire_state_mc_reg_w_lg_q31w(0) AND state_mc_reg(1));
	write_word_64_67_data_valid <= (wire_write_addr_cntr_w_lg_w_q_range541w564w(0) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_68_6B_data_valid <= (wire_write_addr_cntr_w_lg_w_q_range541w564w(0) AND wire_write_addr_cntr_q(0));
	write_word_7c_7f_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_q(1)) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_7c_7f_inv_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_q(1)) AND wire_write_addr_cntr_q(0));
	write_word_done <= (dprio_pulse AND ((write_word_68_6B_data_valid AND rx_reconfig) OR wire_w_lg_write_word_7c_7f_inv_data_valid551w(0)));
	write_word_preemp1t_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_w_lg_w_q_range547w556w(0)) AND wire_write_addr_cntr_q(0));
	write_word_preemp1ta_data_valid <= '0';
	write_word_preemp1tb_data_valid <= '0';
	write_word_vodctrl_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_w_lg_w_q_range547w556w(0)) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_vodctrla_data_valid <= '0';
	wire_w_cal_channel_address_range129w(0) <= cal_channel_address(0);
	wire_w_cal_channel_address_range113w(0) <= cal_channel_address(1);
	wire_w_cal_channel_address_range98w(0) <= cal_channel_address(2);
	wire_w_cal_quad_address_range189w(0) <= cal_quad_address(0);
	wire_w_channel_address_range122w(0) <= channel_address(0);
	wire_w_channel_address_range107w(0) <= channel_address(1);
	wire_w_logical_pll_sel_num_range119w(0) <= logical_pll_sel_num(0);
	wire_w_logical_pll_sel_num_range103w(0) <= logical_pll_sel_num(1);
	wire_w_reconfig_mode_sel_range76w(0) <= reconfig_mode_sel(0);
	wire_w_reconfig_mode_sel_range78w(0) <= reconfig_mode_sel(1);
	wire_w_reconfig_mode_sel_range81w(0) <= reconfig_mode_sel(2);
	wire_w_rx_eqctrl_range458w(0) <= rx_eqctrl(0);
	wire_w_rx_eqctrl_range451w(0) <= rx_eqctrl(1);
	wire_w_rx_eqctrl_range453w(0) <= rx_eqctrl(2);
	wire_w_rx_eqctrl_range455w(0) <= rx_eqctrl(3);
	wire_w_rx_eqdcgain_range432w(0) <= rx_eqdcgain(0);
	wire_w_rx_eqdcgain_range433w(0) <= rx_eqdcgain(1);
	wire_w_rx_eqdcgain_range429w(0) <= rx_eqdcgain(2);
	wire_w_tx_preemp_0t_range2w(0) <= tx_preemp_0t(4);
	wire_w_tx_preemp_0t_wire_range507w <= tx_preemp_0t_wire(3 DOWNTO 0);
	wire_w_tx_preemp_2t_range4w(0) <= tx_preemp_2t(4);
	wire_w_tx_preemp_2t_wire_range511w <= tx_preemp_2t_wire(3 DOWNTO 0);
	wire_w_tx_vodctrl_range374w(0) <= tx_vodctrl(0);
	wire_w_tx_vodctrl_range371w(0) <= tx_vodctrl(1);
	wire_w_tx_vodctrl_range372w(0) <= tx_vodctrl(2);
	wire_w_w_rx_eqv572w_range623w(0) <= w_rx_eqv572w(0);
	wire_w_w_rx_eqv572w_range624w(0) <= w_rx_eqv572w(1);
	wire_w_w_rx_eqv572w_range627w(0) <= w_rx_eqv572w(2);
	loop44 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy171w175w(i) <= wire_calibration_w_lg_busy171w(0) AND a2gr_dprio_addr(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy171w172w(i) <= wire_calibration_w_lg_busy171w(0) AND a2gr_dprio_data(i);
	END GENERATE loop45;
	wire_calibration_w_lg_w_lg_busy171w178w(0) <= wire_calibration_w_lg_busy171w(0) AND a2gr_dprio_rden;
	wire_calibration_w_lg_w_lg_busy171w181w(0) <= wire_calibration_w_lg_busy171w(0) AND a2gr_dprio_wren;
	wire_calibration_w_lg_w_lg_busy171w184w(0) <= wire_calibration_w_lg_busy171w(0) AND a2gr_dprio_wren_data;
	loop46 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy176w(i) <= wire_calibration_busy AND cal_dprio_address(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy173w(i) <= wire_calibration_busy AND wire_calibration_dprio_dataout(i);
	END GENERATE loop47;
	wire_calibration_w_lg_busy171w(0) <= NOT wire_calibration_busy;
	wire_calibration_reset <= wire_w_lg_offset_cancellation_reset152w(0);
	wire_w_lg_offset_cancellation_reset152w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration :  alt_cal
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 3,
		NUMBER_OF_CHANNELS => 8,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_dprio_dataout,
		dprio_rden => wire_calibration_dprio_rden,
		dprio_wren => wire_calibration_dprio_wren,
		quad_addr => wire_calibration_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_reset,
		retain_addr => wire_calibration_retain_addr,
		start => start,
		testbuses => cal_testbuses,
		transceiver_init => transceiver_init
	  );
	wire_dprio_w_lg_w_lg_w_dataout_range704w705w717w(0) <= wire_dprio_w_lg_w_dataout_range704w705w(0) AND wire_dprio_w_dataout_range707w(0);
	wire_dprio_w_lg_w_dataout_range704w713w(0) <= wire_dprio_w_dataout_range704w(0) AND wire_dprio_w_lg_w_dataout_range707w712w(0);
	wire_dprio_w_lg_w_dataout_range704w708w(0) <= wire_dprio_w_dataout_range704w(0) AND wire_dprio_w_dataout_range707w(0);
	wire_dprio_w_lg_w_dataout_range497w706w(0) <= wire_dprio_w_dataout_range497w(0) AND wire_dprio_w_lg_w_dataout_range704w705w(0);
	wire_dprio_w_lg_w_dataout_range497w716w(0) <= wire_dprio_w_dataout_range497w(0) AND wire_dprio_w_dataout_range704w(0);
	wire_dprio_w_lg_w_dataout_range688w689w(0) <= wire_dprio_w_dataout_range688w(0) AND wire_dprio_w_lg_w_dataout_range684w687w(0);
	wire_dprio_w_lg_busy199w(0) <= NOT wire_dprio_busy;
	wire_dprio_w_lg_w_dataout_range684w687w(0) <= NOT wire_dprio_w_dataout_range684w(0);
	wire_dprio_w_lg_w_dataout_range707w712w(0) <= NOT wire_dprio_w_dataout_range707w(0);
	wire_dprio_w_lg_w_dataout_range704w705w(0) <= NOT wire_dprio_w_dataout_range704w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_dataout_range704w705w717w718w(0) <= wire_dprio_w_lg_w_lg_w_dataout_range704w705w717w(0) OR wire_dprio_w_lg_w_dataout_range497w716w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range704w713w714w(0) <= wire_dprio_w_lg_w_dataout_range704w713w(0) OR wire_dprio_w_lg_w_dataout_range497w706w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range704w708w709w(0) <= wire_dprio_w_lg_w_dataout_range704w708w(0) OR wire_dprio_w_lg_w_dataout_range497w706w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_dataout_range692w693w694w695w(0) <= wire_dprio_w_lg_w_lg_w_dataout_range692w693w694w(0) XOR wire_dprio_w_dataout_range684w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range692w693w694w(0) <= wire_dprio_w_lg_w_dataout_range692w693w(0) XOR wire_dprio_w_dataout_range691w(0);
	wire_dprio_w_lg_w_dataout_range692w693w(0) <= wire_dprio_w_dataout_range692w(0) XOR wire_dprio_w_dataout_range688w(0);
	wire_dprio_address <= wire_calibration_w_lg_w_lg_busy176w177w;
	loop48 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy176w177w(i) <= wire_calibration_w_lg_busy176w(i) OR wire_calibration_w_lg_w_lg_busy171w175w(i);
	END GENERATE loop48;
	wire_dprio_datain <= wire_calibration_w_lg_w_lg_busy173w174w;
	loop49 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy173w174w(i) <= wire_calibration_w_lg_busy173w(i) OR wire_calibration_w_lg_w_lg_busy171w172w(i);
	END GENERATE loop49;
	wire_dprio_rden <= wire_calibration_w_lg_w_lg_busy179w180w(0);
	wire_calibration_w_lg_w_lg_busy179w180w(0) <= (wire_calibration_busy AND wire_calibration_dprio_rden) OR wire_calibration_w_lg_w_lg_busy171w178w(0);
	wire_dprio_wren <= wire_calibration_w_lg_w_lg_busy182w183w(0);
	wire_calibration_w_lg_w_lg_busy182w183w(0) <= (wire_calibration_busy AND wire_calibration_dprio_wren) OR wire_calibration_w_lg_w_lg_busy171w181w(0);
	wire_dprio_wren_data <= wire_calibration_w_lg_w_lg_busy185w186w(0);
	wire_calibration_w_lg_w_lg_busy185w186w(0) <= (wire_calibration_busy AND wire_calibration_retain_addr) OR wire_calibration_w_lg_w_lg_busy171w184w(0);
	wire_dprio_w_dataout_range684w(0) <= wire_dprio_dataout(10);
	wire_dprio_w_dataout_range707w(0) <= wire_dprio_dataout(13);
	wire_dprio_w_dataout_range704w(0) <= wire_dprio_dataout(14);
	wire_dprio_w_dataout_range410w <= wire_dprio_dataout(15 DOWNTO 11);
	wire_dprio_w_dataout_range497w(0) <= wire_dprio_dataout(15);
	wire_dprio_w_dataout_range730w <= wire_dprio_dataout(3 DOWNTO 0);
	wire_dprio_w_dataout_range749w(0) <= wire_dprio_dataout(4);
	wire_dprio_w_dataout_range742w <= wire_dprio_dataout(7 DOWNTO 4);
	wire_dprio_w_dataout_range692w(0) <= wire_dprio_dataout(7);
	wire_dprio_w_dataout_range688w(0) <= wire_dprio_dataout(8);
	wire_dprio_w_dataout_range691w(0) <= wire_dprio_dataout(9);
	wire_dprio_w_dataout_range759w(0) <= wire_dprio_dataout(3);
	dprio :  altpcie_reconfig_4sgx_alt_dprio_2vj
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => wire_dprioout_mux_result(0),
		quad_address => quad_address_out,
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		wren => wire_dprio_wren,
		wren_data => wire_dprio_wren_data
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= ( wire_w_lg_w_lg_cal_busy91w92w & wire_w_lg_w_lg_cal_busy99w100w & wire_w_lg_w_lg_cal_busy114w115w & wire_w_lg_w_lg_cal_busy130w131w);
		END IF;
	END PROCESS;
	wire_address_pres_reg_w_lg_w_lg_w_q_range136w137w138w(0) <= wire_address_pres_reg_w_lg_w_q_range136w137w(0) AND wire_address_pres_reg_w_q_range134w(0);
	loop50 : FOR i IN 0 TO 1 GENERATE 
		wire_address_pres_reg_w_lg_w_q_range140w141w(i) <= wire_address_pres_reg_w_q_range140w(i) AND wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range136w137w138w139w(0);
	END GENERATE loop50;
	wire_address_pres_reg_w_lg_w_q_range136w137w(0) <= wire_address_pres_reg_w_q_range136w(0) AND wire_address_pres_reg_w_q_range135w(0);
	wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range136w137w138w139w(0) <= NOT wire_address_pres_reg_w_lg_w_lg_w_q_range136w137w138w(0);
	wire_address_pres_reg_w_q_range134w(0) <= address_pres_reg(0);
	wire_address_pres_reg_w_q_range140w <= address_pres_reg(1 DOWNTO 0);
	wire_address_pres_reg_w_q_range135w(0) <= address_pres_reg(1);
	wire_address_pres_reg_w_q_range136w(0) <= address_pres_reg(2);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN data_valid_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_data_valid_reg_ena = '1') THEN data_valid_reg <= (NOT (is_illegal_reg_out OR reset_system));
			END IF;
		END IF;
	END PROCESS;
	wire_data_valid_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_pulse_reg_ena = '1') THEN dprio_pulse_reg <= wire_dprio_busy;
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_pulse_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN reconf_mode_sel_reg <= reconfig_mode_sel;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(0) = '1') THEN rx_eqctrl_reg(0) <= wire_rx_eqctrl_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(1) = '1') THEN rx_eqctrl_reg(1) <= wire_rx_eqctrl_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(2) = '1') THEN rx_eqctrl_reg(2) <= wire_rx_eqctrl_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(3) = '1') THEN rx_eqctrl_reg(3) <= wire_rx_eqctrl_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_rx_eqctrl_reg_d <= wire_w_lg_w_lg_read_state681w682w;
	loop51 : FOR i IN 0 TO 3 GENERATE
		wire_rx_eqctrl_reg_ena(i) <= wire_w_lg_w_lg_read_word_68_6B_data_valid678w679w(0);
	END GENERATE loop51;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(0) = '1') THEN rx_equalizer_dcgain_reg(0) <= wire_rx_equalizer_dcgain_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(1) = '1') THEN rx_equalizer_dcgain_reg(1) <= wire_rx_equalizer_dcgain_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(2) = '1') THEN rx_equalizer_dcgain_reg(2) <= wire_rx_equalizer_dcgain_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	wire_rx_equalizer_dcgain_reg_d <= wire_w_lg_w_lg_read_state701w702w;
	loop52 : FOR i IN 0 TO 2 GENERATE
		wire_rx_equalizer_dcgain_reg_ena(i) <= wire_w_lg_w_lg_read_word_64_67_data_valid698w699w(0);
	END GENERATE loop52;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN state_mc_reg <= state_mc_reg_in;
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_lg_q31w(0) <= NOT state_mc_reg(0);
	wire_state_mc_reg_w_lg_q29w(0) <= NOT state_mc_reg(1);
	wire_state_mc_reg_w_q_range55w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range67w(0) <= state_mc_reg(1);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemp_0t_inv_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemp_0t_inv_reg_ena = "1") THEN tx_preemp_0t_inv_reg(0) <= (wire_w_lg_read_state750w(0) OR wire_w_lg_write_state748w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemp_0t_inv_reg_ena(0) <= ((read_word_7c_7f_inv_data_valid AND read_state) OR (write_state AND write_word_7c_7f_inv_data_valid));
	wire_tx_preemp_0t_inv_reg_w_lg_w_q_range752w753w(0) <= NOT wire_tx_preemp_0t_inv_reg_w_q_range752w(0);
	wire_tx_preemp_0t_inv_reg_w_q_range752w(0) <= tx_preemp_0t_inv_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemp_2t_inv_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemp_2t_inv_reg_ena = "1") THEN tx_preemp_2t_inv_reg(0) <= (wire_w_lg_read_state760w(0) OR wire_w_lg_write_state758w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemp_2t_inv_reg_ena(0) <= ((read_word_7c_7f_inv_data_valid AND read_state) OR (write_state AND write_word_7c_7f_inv_data_valid));
	wire_tx_preemp_2t_inv_reg_w_lg_w_q_range762w763w(0) <= NOT wire_tx_preemp_2t_inv_reg_w_q_range762w(0);
	wire_tx_preemp_2t_inv_reg_w_q_range762w(0) <= tx_preemp_2t_inv_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(0) = '1') THEN tx_preemphasisctrl_1stposttap_reg(0) <= wire_tx_preemphasisctrl_1stposttap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(1) = '1') THEN tx_preemphasisctrl_1stposttap_reg(1) <= wire_tx_preemphasisctrl_1stposttap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(2) = '1') THEN tx_preemphasisctrl_1stposttap_reg(2) <= wire_tx_preemphasisctrl_1stposttap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(3) = '1') THEN tx_preemphasisctrl_1stposttap_reg(3) <= wire_tx_preemphasisctrl_1stposttap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(4) = '1') THEN tx_preemphasisctrl_1stposttap_reg(4) <= wire_tx_preemphasisctrl_1stposttap_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_1stposttap_reg_d <= wire_w_lg_w_lg_read_state737w738w;
	loop53 : FOR i IN 0 TO 4 GENERATE
		wire_tx_preemphasisctrl_1stposttap_reg_ena(i) <= wire_w_lg_w_lg_read_word_preemp_1t_data_valid734w735w(0);
	END GENERATE loop53;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(0) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(0) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(1) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(1) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(2) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(2) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(3) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(3) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_2ndposttap_reg_d <= wire_w_lg_w_lg_read_state743w744w;
	loop54 : FOR i IN 0 TO 3 GENERATE
		wire_tx_preemphasisctrl_2ndposttap_reg_ena(i) <= wire_w_lg_w_lg_read_word_7c_7f_data_valid739w740w(0);
	END GENERATE loop54;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(0) = '1') THEN tx_preemphasisctrl_pretap_reg(0) <= wire_tx_preemphasisctrl_pretap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(1) = '1') THEN tx_preemphasisctrl_pretap_reg(1) <= wire_tx_preemphasisctrl_pretap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(2) = '1') THEN tx_preemphasisctrl_pretap_reg(2) <= wire_tx_preemphasisctrl_pretap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(3) = '1') THEN tx_preemphasisctrl_pretap_reg(3) <= wire_tx_preemphasisctrl_pretap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_pretap_reg_d <= wire_w_lg_w_lg_read_state731w732w;
	loop55 : FOR i IN 0 TO 3 GENERATE
		wire_tx_preemphasisctrl_pretap_reg_ena(i) <= wire_w_lg_w_lg_read_state727w728w(0);
	END GENERATE loop55;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(0) = '1') THEN tx_vodctrl_reg(0) <= wire_tx_vodctrl_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(1) = '1') THEN tx_vodctrl_reg(1) <= wire_tx_vodctrl_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(2) = '1') THEN tx_vodctrl_reg(2) <= wire_tx_vodctrl_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_vodctrl_reg_d <= wire_w_lg_w_lg_read_state724w725w;
	loop56 : FOR i IN 0 TO 2 GENERATE
		wire_tx_vodctrl_reg_ena(i) <= wire_w_lg_w_lg_read_word_vodctrl_data_valid721w722w(0);
	END GENERATE loop56;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_addr_inc_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN wr_addr_inc_reg <= (wr_pulse OR ((wire_w_lg_wr_pulse144w(0) AND wire_w_lg_rd_pulse143w(0)) AND wr_addr_inc_reg));
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_rd_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wr_rd_pulse_reg_ena = '1') THEN 
				IF (wire_wr_rd_pulse_reg_sclr = '1') THEN wr_rd_pulse_reg <= '0';
				ELSE wr_rd_pulse_reg <= wire_wr_rd_pulse_reg_w_lg_q202w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_wr_rd_pulse_reg_ena <= (dprio_pulse AND wire_w_lg_read_state203w(0));
	wire_wr_rd_pulse_reg_sclr <= (((wire_w_lg_reset_system207w(0) OR (is_diff_mif AND write_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_w_lg_q250w(0) <= wr_rd_pulse_reg AND wire_w_lg_w_lg_is_tier_1222w249w(0);
	wire_wr_rd_pulse_reg_w_lg_q202w(0) <= NOT wr_rd_pulse_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wren_data_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wren_data_reg_ena = '1') THEN wren_data_reg <= (wire_wren_data_reg_w_lg_w_lg_q337w338w(0) OR wire_wren_data_reg_w_lg_q336w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_wren_data_reg_ena <= (is_tier_1 AND (wire_w_lg_is_diff_mif196w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	wire_wren_data_reg_w_lg_w_lg_q337w338w(0) <= wire_wren_data_reg_w_lg_q337w(0) AND rd_pulse;
	wire_wren_data_reg_w_lg_q336w(0) <= wren_data_reg AND wire_w_lg_write_done229w(0);
	wire_wren_data_reg_w_lg_q337w(0) <= NOT wren_data_reg;
	wire_wren_data_reg_w_lg_q341w(0) <= wren_data_reg OR is_analog_control;
	wire_add_sub1_dataa <= (OTHERS => '0');
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => tx_preemp_0t(4),
		dataa => wire_add_sub1_dataa,
		datab => tx_preemp_0t(3 DOWNTO 0),
		result => wire_add_sub1_result
	  );
	wire_add_sub10_add_sub <= wire_tx_preemp_0t_inv_reg_w_lg_w_q_range752w753w(0);
	wire_add_sub10_dataa <= (OTHERS => '0');
	add_sub10 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => wire_add_sub10_add_sub,
		dataa => wire_add_sub10_dataa,
		datab => tx_preemp_0t_out_wire(3 DOWNTO 0),
		result => wire_add_sub10_result
	  );
	wire_add_sub11_add_sub <= wire_tx_preemp_2t_inv_reg_w_lg_w_q_range762w763w(0);
	wire_add_sub11_dataa <= (OTHERS => '0');
	add_sub11 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => wire_add_sub11_add_sub,
		dataa => wire_add_sub11_dataa,
		datab => tx_preemp_2t_out_wire(3 DOWNTO 0),
		result => wire_add_sub11_result
	  );
	wire_add_sub2_dataa <= (OTHERS => '0');
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => tx_preemp_2t(4),
		dataa => wire_add_sub2_dataa,
		datab => tx_preemp_2t(3 DOWNTO 0),
		result => wire_add_sub2_result
	  );
	wire_cmpr6_datab <= "1010";
	cmpr6 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr6_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr6_datab
	  );
	wire_cmpr7_datab <= "0110";
	cmpr7 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr7_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr7_datab
	  );
	wire_cmpr8_datab <= "0011";
	cmpr8 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr8_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr8_datab
	  );
	wire_cmpr9_datab <= (OTHERS => '0');
	cmpr9 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr9_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr9_datab
	  );
	wire_addr_cntr_sclr <= wire_w_lg_write_done256w(0);
	wire_w_lg_write_done256w(0) <= write_done OR reconfig_reset_all;
	wire_addr_cntr_sload <= wire_w_lg_idle_state258w(0);
	wire_w_lg_idle_state258w(0) <= idle_state AND (write_all OR read);
	addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 8,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 3
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_gnd,
		data => logical_channel_address,
		q => wire_addr_cntr_q,
		sclr => wire_addr_cntr_sclr,
		sload => wire_addr_cntr_sload
	  );
	wire_read_addr_cntr_w_lg_w_q_range307w310w(0) <= wire_read_addr_cntr_w_q_range307w(0) AND wire_read_addr_cntr_w_q_range305w(0);
	wire_read_addr_cntr_w_lg_w_q_range305w308w(0) <= wire_read_addr_cntr_w_q_range305w(0) AND wire_read_addr_cntr_w_q_range307w(0);
	wire_read_addr_cntr_w_lg_w_q_range305w321w(0) <= NOT wire_read_addr_cntr_w_q_range305w(0);
	wire_read_addr_cntr_w_lg_w_q_range311w312w(0) <= wire_read_addr_cntr_w_q_range311w(0) OR wire_read_addr_cntr_w_lg_w_q_range307w310w(0);
	wire_read_addr_cntr_cnt_en <= wire_w_lg_read_addr_inc285w(0);
	wire_w_lg_read_addr_inc285w(0) <= read_addr_inc AND is_analog_control;
	wire_read_addr_cntr_data <= ( wire_w_lg_tx_reconfig294w & "0" & "0");
	wire_read_addr_cntr_sclr <= wire_w_lg_w_lg_read_done286w287w(0);
	wire_w_lg_w_lg_read_done286w287w(0) <= (read_done OR reset_system) OR reconfig_reset_all;
	wire_read_addr_cntr_sload <= wire_w_lg_w_lg_idle_state295w296w(0);
	wire_w_lg_w_lg_idle_state295w296w(0) <= (idle_state AND read) AND wire_w_lg_tx_reconfig294w(0);
	wire_read_addr_cntr_w_q_range307w(0) <= wire_read_addr_cntr_q(0);
	wire_read_addr_cntr_w_q_range311w(0) <= wire_read_addr_cntr_q(1);
	wire_read_addr_cntr_w_q_range305w(0) <= wire_read_addr_cntr_q(2);
	read_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 6,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 3
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_read_addr_cntr_cnt_en,
		data => wire_read_addr_cntr_data,
		q => wire_read_addr_cntr_q,
		sclr => wire_read_addr_cntr_sclr,
		sload => wire_read_addr_cntr_sload
	  );
	wire_write_addr_cntr_w_lg_w_q_range543w546w(0) <= wire_write_addr_cntr_w_q_range543w(0) AND wire_write_addr_cntr_w_q_range541w(0);
	wire_write_addr_cntr_w_lg_w_q_range541w564w(0) <= wire_write_addr_cntr_w_q_range541w(0) AND wire_write_addr_cntr_w_lg_w_q_range547w556w(0);
	wire_write_addr_cntr_w_lg_w_q_range541w544w(0) <= wire_write_addr_cntr_w_q_range541w(0) AND wire_write_addr_cntr_w_q_range543w(0);
	wire_write_addr_cntr_w_lg_w_q_range547w556w(0) <= NOT wire_write_addr_cntr_w_q_range547w(0);
	wire_write_addr_cntr_w_lg_w_q_range547w548w(0) <= wire_write_addr_cntr_w_q_range547w(0) OR wire_write_addr_cntr_w_lg_w_q_range543w546w(0);
	wire_write_addr_cntr_data <= ( wire_w_lg_tx_reconfig294w & "0" & "0");
	wire_write_addr_cntr_sclr <= wire_w_lg_w_lg_write_done523w524w(0);
	wire_w_lg_w_lg_write_done523w524w(0) <= (write_done OR reset_system) OR reconfig_reset_all;
	wire_write_addr_cntr_sload <= wire_w_lg_w_lg_idle_state531w532w(0);
	wire_w_lg_w_lg_idle_state531w532w(0) <= (idle_state AND write_all) AND wire_w_lg_tx_reconfig294w(0);
	wire_write_addr_cntr_w_q_range543w(0) <= wire_write_addr_cntr_q(0);
	wire_write_addr_cntr_w_q_range547w(0) <= wire_write_addr_cntr_q(1);
	wire_write_addr_cntr_w_q_range541w(0) <= wire_write_addr_cntr_q(2);
	write_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 6,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 3
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => write_addr_inc,
		data => wire_write_addr_cntr_data,
		q => wire_write_addr_cntr_q,
		sclr => wire_write_addr_cntr_sclr,
		sload => wire_write_addr_cntr_sload
	  );
	chl_addr_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => wire_addr_cntr_q,
		eq => wire_chl_addr_decode_eq
	  );
	reconf_mode_dec :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => reconf_mode_sel_reg,
		eq => wire_reconf_mode_dec_eq
	  );
	aeq_ch_done_mux :  altpcie_reconfig_4sgx_mux_c6a
	  PORT MAP ( 
		data => aeq_ch_done,
		result => wire_aeq_ch_done_mux_result,
		sel => w334w(2 DOWNTO 0)
	  );
	wire_dprioout_mux_sel <= wire_w_lg_w_lg_cal_busy190w191w;
	wire_w_lg_w_lg_cal_busy190w191w(0) <= wire_w_lg_cal_busy190w(0) OR (wire_w_lg_cal_busy89w(0) AND quad_address(0));
	dprioout_mux :  altpcie_reconfig_4sgx_mux_46a
	  PORT MAP ( 
		data => cal_dprioout_wire,
		result => wire_dprioout_mux_result,
		sel => wire_dprioout_mux_sel
	  );

 END RTL; --altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altpcie_reconfig_4sgx IS
	PORT
	(
		logical_channel_address		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		offset_cancellation_reset		: IN STD_LOGIC  := '0';
		read		: IN STD_LOGIC ;
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (33 DOWNTO 0);
		rx_eqctrl		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqdcgain		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		tx_preemp_0t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_1t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_2t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_vodctrl		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		write_all		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqctrl_out		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqdcgain_out		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		tx_preemp_0t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_1t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_2t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_vodctrl_out		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END altpcie_reconfig_4sgx;


ARCHITECTURE RTL OF altpcie_reconfig_4sgx IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt2gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "base_port_width=1;cbx_blackbox_list=-lpm_mux;channel_address_width=3;enable_chl_addr_for_analog_ctrl=TRUE;intended_device_family=Stratix IV;number_of_channels=8;number_of_reconfig_ports=2;read_base_port_width=1;rx_eqdcgain_port_width=3;tx_preemp_port_width=5;enable_buf_cal=true;reconfig_fromgxb_width=34;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire9_bv	: BIT_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (2 DOWNTO 0);



	COMPONENT altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1
	PORT (
			logical_channel_address	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_preemp_1t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_preemp_2t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_vodctrl_out	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			data_valid	: OUT STD_LOGIC ;
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (33 DOWNTO 0);
			tx_preemp_2t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_vodctrl	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_clk	: IN STD_LOGIC ;
			tx_preemp_0t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			rx_eqctrl_out	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_preemp_0t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_preemp_1t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			write_all	: IN STD_LOGIC ;
			read	: IN STD_LOGIC ;
			reconfig_mode_sel	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			rx_eqctrl	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_eqdcgain_out	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			offset_cancellation_reset	: IN STD_LOGIC ;
			rx_eqdcgain	: IN STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire9_bv(2 DOWNTO 0) <= "000";
	sub_wire9    <= To_stdlogicvector(sub_wire9_bv);
	reconfig_togxb    <= sub_wire0(3 DOWNTO 0);
	tx_preemp_2t_out    <= sub_wire1(4 DOWNTO 0);
	tx_vodctrl_out    <= sub_wire2(2 DOWNTO 0);
	data_valid    <= sub_wire3;
	tx_preemp_0t_out    <= sub_wire4(4 DOWNTO 0);
	busy    <= sub_wire5;
	rx_eqctrl_out    <= sub_wire6(3 DOWNTO 0);
	tx_preemp_1t_out    <= sub_wire7(4 DOWNTO 0);
	rx_eqdcgain_out    <= sub_wire8(2 DOWNTO 0);

	altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1_component : altpcie_reconfig_4sgx_alt2gxb_reconfig_squ1
	PORT MAP (
		logical_channel_address => logical_channel_address,
		tx_preemp_1t => tx_preemp_1t,
		reconfig_fromgxb => reconfig_fromgxb,
		tx_preemp_2t => tx_preemp_2t,
		tx_vodctrl => tx_vodctrl,
		reconfig_clk => reconfig_clk,
		tx_preemp_0t => tx_preemp_0t,
		write_all => write_all,
		read => read,
		reconfig_mode_sel => sub_wire9,
		rx_eqctrl => rx_eqctrl,
		offset_cancellation_reset => offset_cancellation_reset,
		rx_eqdcgain => rx_eqdcgain,
		reconfig_togxb => sub_wire0,
		tx_preemp_2t_out => sub_wire1,
		tx_vodctrl_out => sub_wire2,
		data_valid => sub_wire3,
		tx_preemp_0t_out => sub_wire4,
		busy => sub_wire5,
		rx_eqctrl_out => sub_wire6,
		tx_preemp_1t_out => sub_wire7,
		rx_eqdcgain_out => sub_wire8
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: PMA NUMERIC "1"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: CHANNEL_ADDRESS_WIDTH NUMERIC "3"
-- Retrieval info: CONSTANT: ENABLE_CHL_ADDR_FOR_ANALOG_CTRL STRING "TRUE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "8"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "2"
-- Retrieval info: CONSTANT: READ_BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RX_EQDCGAIN_PORT_WIDTH NUMERIC "3"
-- Retrieval info: CONSTANT: TX_PREEMP_PORT_WIDTH NUMERIC "5"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "34"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: USED_PORT: logical_channel_address 0 0 3 0 INPUT NODEFVAL "logical_channel_address[2..0]"
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 34 0 INPUT NODEFVAL "reconfig_fromgxb[33..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: rx_eqctrl 0 0 4 0 INPUT NODEFVAL "rx_eqctrl[3..0]"
-- Retrieval info: USED_PORT: rx_eqctrl_out 0 0 4 0 OUTPUT NODEFVAL "rx_eqctrl_out[3..0]"
-- Retrieval info: USED_PORT: rx_eqdcgain 0 0 3 0 INPUT NODEFVAL "rx_eqdcgain[2..0]"
-- Retrieval info: USED_PORT: rx_eqdcgain_out 0 0 3 0 OUTPUT NODEFVAL "rx_eqdcgain_out[2..0]"
-- Retrieval info: USED_PORT: tx_preemp_0t 0 0 5 0 INPUT NODEFVAL "tx_preemp_0t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_0t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_0t_out[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_1t 0 0 5 0 INPUT NODEFVAL "tx_preemp_1t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_1t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_1t_out[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_2t 0 0 5 0 INPUT NODEFVAL "tx_preemp_2t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_2t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_2t_out[4..0]"
-- Retrieval info: USED_PORT: tx_vodctrl 0 0 3 0 INPUT NODEFVAL "tx_vodctrl[2..0]"
-- Retrieval info: USED_PORT: tx_vodctrl_out 0 0 3 0 OUTPUT NODEFVAL "tx_vodctrl_out[2..0]"
-- Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
-- Retrieval info: CONNECT: @logical_channel_address 0 0 3 0 logical_channel_address 0 0 3 0
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 34 0 reconfig_fromgxb 0 0 34 0
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 3 0 GND 0 0 3 0
-- Retrieval info: CONNECT: @rx_eqctrl 0 0 4 0 rx_eqctrl 0 0 4 0
-- Retrieval info: CONNECT: @rx_eqdcgain 0 0 3 0 rx_eqdcgain 0 0 3 0
-- Retrieval info: CONNECT: @tx_preemp_0t 0 0 5 0 tx_preemp_0t 0 0 5 0
-- Retrieval info: CONNECT: @tx_preemp_1t 0 0 5 0 tx_preemp_1t 0 0 5 0
-- Retrieval info: CONNECT: @tx_preemp_2t 0 0 5 0 tx_preemp_2t 0 0 5 0
-- Retrieval info: CONNECT: @tx_vodctrl 0 0 3 0 tx_vodctrl 0 0 3 0
-- Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: rx_eqctrl_out 0 0 4 0 @rx_eqctrl_out 0 0 4 0
-- Retrieval info: CONNECT: rx_eqdcgain_out 0 0 3 0 @rx_eqdcgain_out 0 0 3 0
-- Retrieval info: CONNECT: tx_preemp_0t_out 0 0 5 0 @tx_preemp_0t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_preemp_1t_out 0 0 5 0 @tx_preemp_1t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_preemp_2t_out 0 0 5 0 @tx_preemp_2t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_vodctrl_out 0 0 3 0 @tx_vodctrl_out 0 0 3 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.v TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx_inst.v FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx_bb.v FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_4sgx_inst.vhd FALSE
