-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb_reconfig 

-- ============================================================
-- File Name: altpcie_reconfig_3cgx.vhd
-- Megafunction Name(s):
-- 			alt_c3gxb_reconfig
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Internal Build 134 03/09/2011 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt_c3gxb_reconfig CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV GX" ENABLE_BUF_CAL="TRUE" NUMBER_OF_CHANNELS=4 NUMBER_OF_RECONFIG_PORTS=1 RECONFIG_FROMGXB_WIDTH=5 RECONFIG_TOGXB_WIDTH=4 busy offset_cancellation_reset reconfig_clk reconfig_fromgxb reconfig_togxb
--VERSION_BEGIN 11.0 cbx_alt_c3gxb_reconfig 2011:03:09:22:37:51:SJ cbx_alt_cal 2011:03:09:22:37:51:SJ cbx_alt_dprio 2011:03:09:22:37:51:SJ cbx_altsyncram 2011:03:09:22:37:54:SJ cbx_cycloneii 2011:03:09:22:37:55:SJ cbx_lpm_add_sub 2011:03:09:22:37:56:SJ cbx_lpm_compare 2011:03:09:22:37:56:SJ cbx_lpm_counter 2011:03:09:22:37:56:SJ cbx_lpm_decode 2011:03:09:22:37:56:SJ cbx_lpm_mux 2011:03:09:22:37:56:SJ cbx_lpm_shiftreg 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ cbx_stratix 2011:03:09:22:37:58:SJ cbx_stratixii 2011:03:09:22:37:58:SJ cbx_stratixiii 2011:03:09:22:37:58:SJ cbx_stratixv 2011:03:09:22:37:58:SJ cbx_util_mgl 2011:03:09:22:37:57:SJ  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone IV GX" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset wren wren_data
--VERSION_BEGIN 11.0 cbx_alt_dprio 2011:03:09:22:37:51:SJ cbx_cycloneii 2011:03:09:22:37:55:SJ cbx_lpm_add_sub 2011:03:09:22:37:56:SJ cbx_lpm_compare 2011:03:09:22:37:56:SJ cbx_lpm_counter 2011:03:09:22:37:56:SJ cbx_lpm_decode 2011:03:09:22:37:56:SJ cbx_lpm_shiftreg 2011:03:09:22:37:56:SJ cbx_mgl 2011:03:09:22:48:24:SJ cbx_stratix 2011:03:09:22:37:58:SJ cbx_stratixii 2011:03:09:22:37:58:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_3cgx_alt_dprio_v5k IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END altpcie_reconfig_3cgx_alt_dprio_v5k;

 ARCHITECTURE RTL OF altpcie_reconfig_3cgx_alt_dprio_v5k IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range453w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range457w463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range457w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range449w450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range449w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range449w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range457w458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb210w387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb210w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_049w50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_068w69w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_084w85w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren38w61w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren38w61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state209w213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state389w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_049w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_068w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_084w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren38w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren38w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren38w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden445w446w447w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state209w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden445w446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden36w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden445w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_049w50w51w(0) <= wire_dprio_w_lg_w_lg_s0_to_049w50w(0) AND wire_state_mc_reg_w_q_range47w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_068w69w70w(0) <= wire_dprio_w_lg_w_lg_s1_to_068w69w(0) AND wire_state_mc_reg_w_q_range66w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_084w85w86w(0) <= wire_dprio_w_lg_w_lg_s2_to_084w85w(0) AND wire_state_mc_reg_w_q_range82w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren38w61w74w(0) <= wire_dprio_w_lg_w_lg_wren38w61w(0) AND wire_dprio_w_lg_rdinc73w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren38w61w62w(0) <= wire_dprio_w_lg_w_lg_wren38w61w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state209w213w214w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state209w213w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state389w390w(0) <= wire_dprio_w_lg_rd_data_output_state389w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state324w325w(0) <= wire_dprio_w_lg_wr_data_state324w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_049w50w(0) <= wire_dprio_w_lg_s0_to_049w(0) AND wire_dprio_w_lg_s0_to_148w(0);
	wire_dprio_w_lg_w_lg_s1_to_068w69w(0) <= wire_dprio_w_lg_s1_to_068w(0) AND wire_dprio_w_lg_s1_to_167w(0);
	wire_dprio_w_lg_w_lg_s2_to_084w85w(0) <= wire_dprio_w_lg_s2_to_084w(0) AND wire_dprio_w_lg_s2_to_183w(0);
	wire_dprio_w_lg_w_lg_wren38w61w(0) <= wire_dprio_w_lg_wren38w(0) AND wire_dprio_w_lg_wren_data60w(0);
	wire_dprio_w_lg_w_lg_wren38w39w(0) <= wire_dprio_w_lg_wren38w(0) AND wire_dprio_w_lg_w_lg_rden36w37w(0);
	wire_dprio_w_lg_w_lg_wren38w56w(0) <= wire_dprio_w_lg_wren38w(0) AND wire_dprio_w_lg_rdinc55w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden445w446w447w448w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden445w446w447w(0) AND wire_dprio_w_lg_startup_done443w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state209w213w(0) <= wire_dprio_w_lg_wr_addr_state209w(0) AND wire_addr_shift_reg_w_q_range212w(0);
	wire_dprio_w_lg_idle_state75w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren38w61w74w(0);
	wire_dprio_w_lg_idle_state57w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren38w56w(0);
	wire_dprio_w_lg_idle_state64w(0) <= idle_state AND wire_dprio_w_lg_wren63w(0);
	wire_dprio_w_lg_idle_state41w(0) <= idle_state AND wire_dprio_w_lg_wren40w(0);
	wire_dprio_w_lg_idle_state78w(0) <= idle_state AND wire_dprio_w_lg_wren77w(0);
	wire_dprio_w_lg_rd_data_output_state389w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range388w(0);
	wire_dprio_w_lg_wr_data_state324w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range323w(0);
	wire_dprio_w_lg_s0_to_049w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_148w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_068w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_167w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_084w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_183w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done443w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle444w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren38w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data60w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden445w446w447w(0) <= wire_dprio_w_lg_w_lg_rden445w446w(0) OR wire_dprio_w_lg_startup_idle444w(0);
	wire_dprio_w_lg_w_lg_rden36w37w(0) <= wire_dprio_w_lg_rden36w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden445w446w(0) <= wire_dprio_w_lg_rden445w(0) OR rdinc;
	wire_dprio_w_lg_rden36w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden445w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc73w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc55w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_152w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_049w50w51w(0);
	wire_dprio_w_lg_s1_to_171w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_068w69w70w(0);
	wire_dprio_w_lg_s2_to_187w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_084w85w86w(0);
	wire_dprio_w_lg_wr_addr_state209w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren63w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren38w61w62w(0);
	wire_dprio_w_lg_wren40w(0) <= wren OR wire_dprio_w_lg_w_lg_wren38w39w(0);
	wire_dprio_w_lg_wren77w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range457w466w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range449w454w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state41w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state64w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state57w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state78w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state75w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range457w463w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range449w450w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range212w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range388w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range457w458w & wire_startup_cntr_w_lg_w_q_range449w454w & wire_startup_cntr_w_lg_w_q_range449w450w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden445w446w447w448w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range453w456w(0) <= wire_startup_cntr_w_q_range453w(0) AND wire_startup_cntr_w_q_range449w(0);
	wire_startup_cntr_w_lg_w_q_range457w463w(0) <= wire_startup_cntr_w_q_range457w(0) AND wire_startup_cntr_w_lg_w_q_range449w450w(0);
	wire_startup_cntr_w_lg_w_q_range457w466w(0) <= wire_startup_cntr_w_q_range457w(0) AND wire_startup_cntr_w_lg_w_q_range449w465w(0);
	wire_startup_cntr_w_lg_w_q_range449w450w(0) <= NOT wire_startup_cntr_w_q_range449w(0);
	wire_startup_cntr_w_lg_w_q_range449w465w(0) <= wire_startup_cntr_w_q_range449w(0) OR wire_startup_cntr_w_q_range453w(0);
	wire_startup_cntr_w_lg_w_q_range449w454w(0) <= wire_startup_cntr_w_q_range449w(0) XOR wire_startup_cntr_w_q_range453w(0);
	wire_startup_cntr_w_lg_w_q_range457w458w(0) <= wire_startup_cntr_w_q_range457w(0) XOR wire_startup_cntr_w_lg_w_q_range453w456w(0);
	wire_startup_cntr_w_q_range449w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range453w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range457w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_187w & wire_dprio_w_lg_s1_to_171w & wire_dprio_w_lg_s0_to_152w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range47w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range66w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range82w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range323w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb210w387w(0) <= wire_pre_amble_cmpr_w_lg_agb210w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb210w322w(0) <= wire_pre_amble_cmpr_w_lg_agb210w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb210w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state32w(0);
	wire_dprio_w_lg_write_state32w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state209w213w214w(0) OR (wire_pre_amble_cmpr_w_lg_agb210w(0) AND wire_dprio_w_lg_wr_addr_state209w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state324w325w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb210w322w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state389w390w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb210w387w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --altpcie_reconfig_3cgx_alt_dprio_v5k

 LIBRARY altera_mf;
 USE altera_mf.all;

--synthesis_resources = alt_cal_c3gxb 1 lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 114 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 offset_cancellation_reset	:	IN  STD_LOGIC := '0';
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp;

 ARCHITECTURE RTL OF altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0";

	 SIGNAL  wire_calibration_c3gxb_w_lg_busy8w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy7w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_c3gxb_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_c3gxb_w_lg_busy10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 COMPONENT  alt_cal_c3gxb
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_type	:	STRING := "alt_cal_c3gxb"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  altpcie_reconfig_3cgx_alt_dprio_v5k
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	busy <= cal_busy;
	cal_busy <= wire_calibration_c3gxb_busy;
	cal_dprioout_wire(0) <= ( reconfig_fromgxb(0));
	cal_testbuses <= ( reconfig_fromgxb(4 DOWNTO 1));
	channel_address <= wire_calibration_c3gxb_dprio_addr(14 DOWNTO 12);
	dprio_address <= ( wire_calibration_c3gxb_dprio_addr(15) & address_pres_reg(2 DOWNTO 0) & wire_calibration_c3gxb_dprio_addr(11 DOWNTO 0));
	quad_address <= wire_calibration_c3gxb_quad_addr;
	reconfig_reset_all <= '0';
	reconfig_togxb <= ( wire_calibration_c3gxb_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	loop1 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy8w(i) <= wire_calibration_c3gxb_busy AND dprio_address(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_c3gxb_w_lg_busy7w(i) <= wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_dataout(i);
	END GENERATE loop2;
	wire_calibration_c3gxb_reset <= wire_w_lg_offset_cancellation_reset5w(0);
	wire_w_lg_offset_cancellation_reset5w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration_c3gxb :  alt_cal_c3gxb
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 2,
		NUMBER_OF_CHANNELS => 4,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_c3gxb_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_c3gxb_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_c3gxb_dprio_dataout,
		dprio_rden => wire_calibration_c3gxb_dprio_rden,
		dprio_wren => wire_calibration_c3gxb_dprio_wren,
		quad_addr => wire_calibration_c3gxb_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_c3gxb_reset,
		retain_addr => wire_calibration_c3gxb_retain_addr,
		testbuses => cal_testbuses
	  );
	wire_dprio_address <= wire_calibration_c3gxb_w_lg_busy8w;
	wire_dprio_datain <= wire_calibration_c3gxb_w_lg_busy7w;
	wire_dprio_rden <= wire_calibration_c3gxb_w_lg_busy9w(0);
	wire_calibration_c3gxb_w_lg_busy9w(0) <= wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_rden;
	wire_dprio_wren <= wire_calibration_c3gxb_w_lg_busy10w(0);
	wire_calibration_c3gxb_w_lg_busy10w(0) <= wire_calibration_c3gxb_busy AND wire_calibration_c3gxb_dprio_wren;
	dprio :  altpcie_reconfig_3cgx_alt_dprio_v5k
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => cal_dprioout_wire(0),
		quad_address => address_pres_reg(11 DOWNTO 3),
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		wren => wire_dprio_wren,
		wren_data => wire_calibration_c3gxb_retain_addr
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= ( quad_address & channel_address);
		END IF;
	END PROCESS;

 END RTL; --altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altpcie_reconfig_3cgx IS
	PORT
	(
		offset_cancellation_reset		: IN STD_LOGIC  := '0';
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		busy		: OUT STD_LOGIC ;
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END altpcie_reconfig_3cgx;


ARCHITECTURE RTL OF altpcie_reconfig_3cgx IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt_c3gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "cbx_blackbox_list=-lpm_mux;intended_device_family=Cyclone IV GX;number_of_channels=4;number_of_reconfig_ports=1;enable_buf_cal=true;reconfig_fromgxb_width=5;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp
	PORT (
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			offset_cancellation_reset	: IN STD_LOGIC ;
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	reconfig_togxb    <= sub_wire0(3 DOWNTO 0);
	busy    <= sub_wire1;

	altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp_component : altpcie_reconfig_3cgx_alt_c3gxb_reconfig_ffp
	PORT MAP (
		reconfig_clk => reconfig_clk,
		offset_cancellation_reset => offset_cancellation_reset,
		reconfig_fromgxb => reconfig_fromgxb,
		reconfig_togxb => sub_wire0,
		busy => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: PMA NUMERIC "0"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "1"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 INPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 5 0 reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.v TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_inst.v FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_bb.v TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altpcie_reconfig_3cgx_inst.vhd FALSE
