
module clock_buffer (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
